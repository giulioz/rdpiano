module test();

reg [7:0] env_param_5_r;
reg [20:0] adder1_b;

wire adder1_b_high;
assign adder1_b_high = (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7];

initial begin
  env_param_5_r = 8'd0;
  for (integer i = 0; i < 256; i++) begin
    env_param_5_r = i[7:0];
    // env_param_5_r[7:2] = i;
    adder1_b[0] = ~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3] && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[1] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[2] = ~((((~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || ((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~((~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || ((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[3] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[4] = ~((((0 && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || ((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~((0 && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || ((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[5] = ~((~(~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0])) || ~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]))) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || ((~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0])) || ~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]))) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[6] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[7] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[8] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (~env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[9] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[10] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[11] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && ~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[12] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (~env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[13] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[14] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[6] && ~env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[15] = ~(((((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(((~(~env_param_5_r[2] || env_param_5_r[1]) || env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[16] = ~((((((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (0 && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~((((~env_param_5_r[2] && ~env_param_5_r[1] && env_param_5_r[0]) || ~((~env_param_5_r[2] && env_param_5_r[0]) || ~env_param_5_r[1])) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (0 && env_param_5_r[6] && ~env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[17] = ~((((~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~((~(~env_param_5_r[2] && ~env_param_5_r[1]) && ~env_param_5_r[0] && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[18] = ~((((((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~((((env_param_5_r[2] && ~env_param_5_r[1] && ~env_param_5_r[0]) || ~(~env_param_5_r[1] || ~env_param_5_r[0])) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3]) || (env_param_5_r[6] && env_param_5_r[5] && ~env_param_5_r[4] && env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[19] = ~((((env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3])) && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~((env_param_5_r[2] && ~(~env_param_5_r[1] && ~env_param_5_r[0]) && env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) || (env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && ~env_param_5_r[3])) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    adder1_b[20] = ~((env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3] && (env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7]) || (~(env_param_5_r[6] && env_param_5_r[5] && env_param_5_r[4] && env_param_5_r[3]) && ~((env_param_5_r[6] || env_param_5_r[5] || env_param_5_r[4] || env_param_5_r[3]) && (env_param_5_r[2] || env_param_5_r[1] || env_param_5_r[0]) && env_param_5_r[7])));
    $display("%x", adder1_b);
  end
end

endmodule
