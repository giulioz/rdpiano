module cell_1_a();
endmodule
module cell_1_b();
endmodule
module cell_1_c();
endmodule
module cell_1_d();
endmodule
module cell_1_e();
endmodule
module cell_2_a();
endmodule
module cell_2_b();
endmodule
module cell_2_c();
endmodule
module cell_2_d();
endmodule
module cell_2_e();
endmodule
module cell_2_f();
endmodule
module cell_2_g();
endmodule
module cell_2_h();
endmodule
module cell_2_i();
endmodule
module cell_3_a();
endmodule
module cell_3_b();
endmodule
module cell_3_c();
endmodule
module cell_3_d();
endmodule
module cell_3_e();
endmodule
module cell_4_a();
endmodule
module cell_4_b();
endmodule
module cell_4_c();
endmodule
module cell_4_d();
endmodule
module cell_5_a();
endmodule
module cell_6_a();
endmodule
module cell_6_b();
endmodule
module cell_6_c();
endmodule
module cell_6_d();
endmodule
module cell_6_e();
endmodule
module cell_7_a();
endmodule
module cell_7_b();
endmodule
module cell_7_c();
endmodule
module cell_8_fd2_fd7_fdp_a1n_sm1();
endmodule
module cell_9_a();
endmodule
module cell_11_a();
endmodule
module cell_13_lt4();
endmodule
module cell_15_lt3_ltm();
endmodule
module cell_21_fdp();
endmodule
module cell_48_c34_c35();
endmodule
module cell_50_a4h();
endmodule

cell_11_a inst_6_20 ();
cell_13_lt4 inst_0_19 ();
cell_13_lt4 inst_0_3 ();
cell_13_lt4 inst_0_74 ();
cell_13_lt4 inst_10_19 ();
cell_13_lt4 inst_10_2 ();
cell_13_lt4 inst_10_33 ();
cell_13_lt4 inst_13_60 ();
cell_13_lt4 inst_13_76 ();
cell_13_lt4 inst_13_92 ();
cell_13_lt4 inst_14_107 ();
cell_13_lt4 inst_14_60 ();
cell_13_lt4 inst_14_74 ();
cell_13_lt4 inst_14_94 ();
cell_13_lt4 inst_15_91 ();
cell_13_lt4 inst_16_106 ();
cell_13_lt4 inst_17_106 ();
cell_13_lt4 inst_17_60 ();
cell_13_lt4 inst_17_92 ();
cell_13_lt4 inst_18_105 ();
cell_13_lt4 inst_19_16 ();
cell_13_lt4 inst_19_3 ();
cell_13_lt4 inst_19_32 ();
cell_13_lt4 inst_1_60 ();
cell_13_lt4 inst_1_73 ();
cell_13_lt4 inst_1_86 ();
cell_13_lt4 inst_20_30 ();
cell_13_lt4 inst_21_32 ();
cell_13_lt4 inst_21_47 ();
cell_13_lt4 inst_21_60 ();
cell_13_lt4 inst_21_77 ();
cell_15_lt3_ltm inst_13_45 ();
cell_1_a inst_0_2 ();
cell_1_a inst_0_46 ();
cell_1_a inst_0_47 ();
cell_1_a inst_10_15 ();
cell_1_a inst_10_57 ();
cell_1_a inst_12_57 ();
cell_1_a inst_13_14 ();
cell_1_a inst_20_19 ();
cell_1_a inst_20_24 ();
cell_1_a inst_20_29 ();
cell_1_a inst_20_47 ();
cell_1_a inst_20_50 ();
cell_1_a inst_20_53 ();
cell_1_a inst_20_6 ();
cell_1_a inst_20_7 ();
cell_1_a inst_5_91 ();
cell_1_a inst_6_1 ();
cell_1_a inst_6_5 ();
cell_1_a inst_6_62 ();
cell_1_a inst_6_63 ();
cell_1_a inst_6_64 ();
cell_1_a inst_6_65 ();
cell_1_a inst_7_51 ();
cell_1_a inst_7_54 ();
cell_1_a inst_7_55 ();
cell_1_a inst_7_60 ();
cell_1_a inst_7_61 ();
cell_1_a inst_7_62 ();
cell_1_a inst_8_14 ();
cell_1_a inst_8_19 ();
cell_1_a inst_8_27 ();
cell_1_a inst_8_44 ();
cell_1_a inst_8_47 ();
cell_1_a inst_8_48 ();
cell_1_a inst_8_59 ();
cell_1_a inst_9_55 ();
cell_1_b inst_0_17 ();
cell_1_b inst_0_95 ();
cell_1_b inst_10_56 ();
cell_1_b inst_10_60 ();
cell_1_b inst_10_61 ();
cell_1_b inst_10_62 ();
cell_1_b inst_10_63 ();
cell_1_b inst_10_64 ();
cell_1_b inst_10_65 ();
cell_1_b inst_10_81 ();
cell_1_b inst_10_82 ();
cell_1_b inst_10_93 ();
cell_1_b inst_12_52 ();
cell_1_b inst_12_53 ();
cell_1_b inst_12_54 ();
cell_1_b inst_12_55 ();
cell_1_b inst_16_10 ();
cell_1_b inst_16_104 ();
cell_1_b inst_16_119 ();
cell_1_b inst_16_27 ();
cell_1_b inst_16_90 ();
cell_1_b inst_16_91 ();
cell_1_b inst_1_11 ();
cell_1_b inst_20_0 ();
cell_1_b inst_20_11 ();
cell_1_b inst_20_12 ();
cell_1_b inst_20_13 ();
cell_1_b inst_20_14 ();
cell_1_b inst_20_15 ();
cell_1_b inst_20_16 ();
cell_1_b inst_20_43 ();
cell_1_b inst_20_44 ();
cell_1_b inst_20_46 ();
cell_1_b inst_20_60 ();
cell_1_b inst_20_8 ();
cell_1_b inst_20_9 ();
cell_1_b inst_21_0 ();
cell_1_b inst_21_1 ();
cell_1_b inst_21_104 ();
cell_1_b inst_21_119 ();
cell_1_b inst_21_2 ();
cell_1_b inst_21_3 ();
cell_1_b inst_21_30 ();
cell_1_b inst_21_31 ();
cell_1_b inst_21_4 ();
cell_1_b inst_21_45 ();
cell_1_b inst_21_46 ();
cell_1_b inst_21_7 ();
cell_1_b inst_21_73 ();
cell_1_b inst_21_74 ();
cell_1_b inst_21_76 ();
cell_1_b inst_21_8 ();
cell_1_b inst_21_96 ();
cell_1_b inst_21_97 ();
cell_1_b inst_2_0 ();
cell_1_b inst_2_1 ();
cell_1_b inst_2_2 ();
cell_1_b inst_2_68 ();
cell_1_b inst_3_10 ();
cell_1_b inst_3_60 ();
cell_1_b inst_4_113 ();
cell_1_b inst_4_114 ();
cell_1_b inst_4_115 ();
cell_1_b inst_5_5 ();
cell_1_b inst_6_31 ();
cell_1_b inst_6_32 ();
cell_1_b inst_6_33 ();
cell_1_b inst_6_38 ();
cell_1_b inst_6_6 ();
cell_1_b inst_6_7 ();
cell_1_b inst_7_50 ();
cell_1_b inst_7_66 ();
cell_1_b inst_8_46 ();
cell_1_c inst_0_18 ();
cell_1_c inst_0_35 ();
cell_1_c inst_0_38 ();
cell_1_c inst_10_100 ();
cell_1_c inst_10_101 ();
cell_1_c inst_10_102 ();
cell_1_c inst_10_55 ();
cell_1_c inst_10_66 ();
cell_1_c inst_10_95 ();
cell_1_c inst_12_56 ();
cell_1_c inst_14_26 ();
cell_1_c inst_16_1 ();
cell_1_c inst_16_15 ();
cell_1_c inst_16_2 ();
cell_1_c inst_16_5 ();
cell_1_c inst_16_9 ();
cell_1_c inst_19_31 ();
cell_1_c inst_1_8 ();
cell_1_c inst_20_1 ();
cell_1_c inst_20_10 ();
cell_1_c inst_20_17 ();
cell_1_c inst_20_18 ();
cell_1_c inst_20_22 ();
cell_1_c inst_20_23 ();
cell_1_c inst_20_45 ();
cell_1_c inst_21_111 ();
cell_1_c inst_2_9 ();
cell_1_c inst_3_1 ();
cell_1_c inst_3_6 ();
cell_1_c inst_3_61 ();
cell_1_c inst_3_62 ();
cell_1_c inst_3_63 ();
cell_1_c inst_3_7 ();
cell_1_c inst_4_54 ();
cell_1_c inst_4_55 ();
cell_1_c inst_5_2 ();
cell_1_c inst_6_10 ();
cell_1_c inst_6_59 ();
cell_1_c inst_8_26 ();
cell_1_c inst_8_28 ();
cell_1_c inst_8_45 ();
cell_1_d inst_10_104 ();
cell_1_d inst_10_105 ();
cell_1_d inst_10_106 ();
cell_1_d inst_10_107 ();
cell_1_d inst_10_108 ();
cell_1_d inst_10_109 ();
cell_1_d inst_10_77 ();
cell_1_d inst_10_78 ();
cell_1_d inst_10_79 ();
cell_1_d inst_10_80 ();
cell_1_d inst_10_94 ();
cell_1_d inst_10_96 ();
cell_1_d inst_10_97 ();
cell_1_d inst_10_98 ();
cell_1_d inst_10_99 ();
cell_1_d inst_11_19 ();
cell_1_d inst_11_39 ();
cell_1_d inst_11_59 ();
cell_1_d inst_16_28 ();
cell_1_d inst_16_44 ();
cell_1_d inst_16_8 ();
cell_1_d inst_17_119 ();
cell_1_d inst_19_60 ();
cell_1_d inst_19_61 ();
cell_1_d inst_19_62 ();
cell_1_d inst_19_63 ();
cell_1_d inst_19_64 ();
cell_1_d inst_19_65 ();
cell_1_d inst_19_66 ();
cell_1_d inst_21_112 ();
cell_1_d inst_6_2 ();
cell_1_e inst_6_19 ();
cell_21_fdp inst_0_97 ();
cell_21_fdp inst_18_9 ();
cell_21_fdp inst_1_99 ();
cell_21_fdp inst_21_9 ();
cell_21_fdp inst_3_65 ();
cell_21_fdp inst_3_95 ();
cell_21_fdp inst_5_60 ();
cell_21_fdp inst_5_93 ();
cell_2_a inst_0_33 ();
cell_2_a inst_0_36 ();
cell_2_a inst_0_48 ();
cell_2_a inst_0_50 ();
cell_2_a inst_0_52 ();
cell_2_a inst_0_54 ();
cell_2_a inst_0_56 ();
cell_2_a inst_0_58 ();
cell_2_a inst_0_60 ();
cell_2_a inst_0_62 ();
cell_2_a inst_0_64 ();
cell_2_a inst_0_66 ();
cell_2_a inst_0_89 ();
cell_2_a inst_0_91 ();
cell_2_a inst_0_93 ();
cell_2_a inst_10_17 ();
cell_2_a inst_10_58 ();
cell_2_a inst_10_67 ();
cell_2_a inst_10_69 ();
cell_2_a inst_10_71 ();
cell_2_a inst_10_73 ();
cell_2_a inst_11_106 ();
cell_2_a inst_11_108 ();
cell_2_a inst_11_110 ();
cell_2_a inst_11_112 ();
cell_2_a inst_11_93 ();
cell_2_a inst_11_95 ();
cell_2_a inst_11_97 ();
cell_2_a inst_12_100 ();
cell_2_a inst_12_102 ();
cell_2_a inst_12_107 ();
cell_2_a inst_12_109 ();
cell_2_a inst_12_111 ();
cell_2_a inst_12_58 ();
cell_2_a inst_13_12 ();
cell_2_a inst_15_60 ();
cell_2_a inst_15_76 ();
cell_2_a inst_15_78 ();
cell_2_a inst_15_86 ();
cell_2_a inst_15_88 ();
cell_2_a inst_16_60 ();
cell_2_a inst_16_68 ();
cell_2_a inst_16_70 ();
cell_2_a inst_16_72 ();
cell_2_a inst_16_87 ();
cell_2_a inst_17_25 ();
cell_2_a inst_17_87 ();
cell_2_a inst_17_89 ();
cell_2_a inst_18_118 ();
cell_2_a inst_18_80 ();
cell_2_a inst_18_82 ();
cell_2_a inst_18_90 ();
cell_2_a inst_20_2 ();
cell_2_a inst_20_20 ();
cell_2_a inst_20_25 ();
cell_2_a inst_20_27 ();
cell_2_a inst_20_4 ();
cell_2_a inst_20_48 ();
cell_2_a inst_20_51 ();
cell_2_a inst_20_54 ();
cell_2_a inst_2_60 ();
cell_2_a inst_2_62 ();
cell_2_a inst_2_64 ();
cell_2_a inst_2_66 ();
cell_2_a inst_6_3 ();
cell_2_a inst_6_60 ();
cell_2_a inst_7_52 ();
cell_2_a inst_7_56 ();
cell_2_a inst_7_58 ();
cell_2_a inst_7_63 ();
cell_2_a inst_8_114 ();
cell_2_a inst_8_116 ();
cell_2_a inst_8_118 ();
cell_2_a inst_8_15 ();
cell_2_a inst_8_17 ();
cell_2_a inst_8_49 ();
cell_2_a inst_9_56 ();
cell_2_a inst_9_58 ();
cell_2_a inst_9_60 ();
cell_2_a inst_9_62 ();
cell_2_b inst_19_29 ();
cell_2_b inst_1_6 ();
cell_2_b inst_21_109 ();
cell_2_b inst_3_8 ();
cell_2_c inst_14_22 ();
cell_2_c inst_14_24 ();
cell_2_c inst_14_46 ();
cell_2_c inst_16_25 ();
cell_2_c inst_16_3 ();
cell_2_c inst_16_31 ();
cell_2_c inst_19_1 ();
cell_2_c inst_1_9 ();
cell_2_c inst_21_5 ();
cell_2_c inst_2_10 ();
cell_2_c inst_4_116 ();
cell_2_c inst_4_118 ();
cell_2_c inst_5_0 ();
cell_2_c inst_6_34 ();
cell_2_c inst_6_36 ();
cell_2_c inst_6_8 ();
cell_2_d inst_3_2 ();
cell_2_d inst_3_4 ();
cell_2_d inst_4_56 ();
cell_2_e inst_13_15 ();
cell_2_e inst_13_17 ();
cell_2_e inst_13_19 ();
cell_2_e inst_13_21 ();
cell_2_e inst_13_23 ();
cell_2_e inst_13_31 ();
cell_2_e inst_13_33 ();
cell_2_e inst_13_35 ();
cell_2_e inst_13_37 ();
cell_2_e inst_13_39 ();
cell_2_e inst_13_41 ();
cell_2_e inst_13_43 ();
cell_2_e inst_14_48 ();
cell_2_e inst_14_50 ();
cell_2_e inst_14_52 ();
cell_2_e inst_14_54 ();
cell_2_e inst_14_56 ();
cell_2_e inst_14_58 ();
cell_2_e inst_16_6 ();
cell_2_e inst_19_45 ();
cell_2_e inst_21_117 ();
cell_2_e inst_4_58 ();
cell_2_e inst_5_3 ();
cell_2_f inst_5_89 ();
cell_2_f inst_8_57 ();
cell_2_g inst_15_43 ();
cell_2_h inst_16_11 ();
cell_2_h inst_16_33 ();
cell_2_i inst_16_13 ();
cell_2_i inst_16_29 ();
cell_3_a inst_0_39 ();
cell_3_a inst_0_42 ();
cell_3_b inst_13_1 ();
cell_3_b inst_6_53 ();
cell_3_b inst_6_56 ();
cell_3_c inst_10_110 ();
cell_3_c inst_10_113 ();
cell_3_c inst_10_116 ();
cell_3_c inst_10_83 ();
cell_3_d inst_18_0 ();
cell_3_d inst_18_3 ();
cell_3_d inst_18_30 ();
cell_3_d inst_18_33 ();
cell_3_d inst_18_36 ();
cell_3_d inst_18_39 ();
cell_3_d inst_18_42 ();
cell_3_d inst_18_45 ();
cell_3_d inst_18_48 ();
cell_3_d inst_18_51 ();
cell_3_d inst_18_54 ();
cell_3_d inst_18_57 ();
cell_3_d inst_18_6 ();
cell_3_d inst_19_47 ();
cell_3_d inst_19_50 ();
cell_3_d inst_19_53 ();
cell_3_e inst_21_106 ();
cell_48_c34_c45 inst_1_12 ();
cell_48_c34_c45 inst_2_12 ();
cell_48_c34_c45 inst_3_12 ();
cell_48_c34_c45 inst_4_6 ();
cell_48_c34_c45 inst_5_12 ();
cell_4_a inst_0_68 ();
cell_4_a inst_10_47 ();
cell_4_a inst_10_51 ();
cell_4_b inst_21_113 ();
cell_4_b inst_3_90 ();
cell_4_b inst_4_1 ();
cell_4_c inst_13_4 ();
cell_4_c inst_13_8 ();
cell_4_c inst_14_10 ();
cell_4_c inst_14_2 ();
cell_4_c inst_14_27 ();
cell_4_c inst_14_6 ();
cell_4_c inst_15_111 ();
cell_4_c inst_15_115 ();
cell_4_c inst_6_45 ();
cell_4_c inst_6_49 ();
cell_4_d inst_19_56 ();
cell_4_d inst_20_56 ();
cell_50_a4h inst_12_2 ();
cell_50_a4h inst_19_68 ();
cell_50_a4h inst_20_68 ();
cell_50_a4h inst_2_70 ();
cell_50_a4h inst_4_60 ();
cell_50_a4h inst_6_67 ();
cell_50_a4h inst_7_0 ();
cell_50_a4h inst_7_68 ();
cell_50_a4h inst_8_60 ();
cell_50_a4h inst_9_5 ();
cell_50_a4h inst_9_65 ();
cell_5_a inst_13_114 ();
cell_6_a inst_10_86 ();
cell_6_a inst_11_114 ();
cell_6_a inst_11_60 ();
cell_6_a inst_11_66 ();
cell_6_a inst_11_74 ();
cell_6_a inst_11_80 ();
cell_6_a inst_11_86 ();
cell_6_a inst_11_99 ();
cell_6_a inst_12_113 ();
cell_6_a inst_12_60 ();
cell_6_a inst_12_66 ();
cell_6_a inst_12_74 ();
cell_6_a inst_12_80 ();
cell_6_a inst_12_88 ();
cell_6_a inst_12_94 ();
cell_6_a inst_15_62 ();
cell_6_a inst_15_68 ();
cell_6_a inst_15_80 ();
cell_6_a inst_16_62 ();
cell_6_a inst_16_75 ();
cell_6_a inst_16_81 ();
cell_6_a inst_16_92 ();
cell_6_a inst_16_98 ();
cell_6_a inst_18_60 ();
cell_6_a inst_18_66 ();
cell_6_a inst_18_72 ();
cell_6_a inst_18_84 ();
cell_6_a inst_18_98 ();
cell_6_a inst_1_0 ();
cell_6_a inst_21_98 ();
cell_6_a inst_2_3 ();
cell_6_a inst_5_6 ();
cell_6_a inst_6_39 ();
cell_6_b inst_13_25 ();
cell_6_b inst_14_32 ();
cell_6_c inst_13_108 ();
cell_6_c inst_14_87 ();
cell_6_c inst_15_105 ();
cell_6_c inst_17_75 ();
cell_6_c inst_17_81 ();
cell_6_c inst_18_92 ();
cell_6_c inst_20_61 ();
cell_6_c inst_21_90 ();
cell_6_d inst_15_45 ();
cell_6_d inst_17_10 ();
cell_6_d inst_17_45 ();
cell_6_e inst_16_45 ();
cell_7_a inst_14_15 ();
cell_7_b inst_14_38 ();
cell_7_c inst_15_27 ();
cell_8_fd2_fd7_fdp_a1n_sm1 inst_6_11 ();
cell_9_a inst_15_0 ();
cell_9_a inst_15_18 ();
cell_9_a inst_15_34 ();
cell_9_a inst_15_51 ();
cell_9_a inst_15_9 ();
cell_9_a inst_16_16 ();
cell_9_a inst_16_35 ();
cell_9_a inst_16_51 ();
cell_9_a inst_17_1 ();
cell_9_a inst_17_16 ();
cell_9_a inst_17_27 ();
cell_9_a inst_17_36 ();
cell_9_a inst_17_51 ();
