module test();

reg [7:0] env_speed_r;
reg [20:0] adder1_b;
reg env_speed_some_high;
reg adder1_b_invert;
reg env_mystery;

initial begin
  env_speed_r = 8'd0;
  for (integer i = 0; i < 256; i++) begin
    env_speed_r = i[7:0];
    // env_speed_r = 8'h80;

    // env_speed_some_high = (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3]) && (env_speed_r[2] || env_speed_r[1] || env_speed_r[0]);
    // adder1_b_invert = env_speed_some_high && env_speed_r[7];
    // adder1_b[0] = !(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3] && adder1_b_invert) || (!((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) && !(adder1_b_invert)));
    // adder1_b[1] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[2] = !((((!env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || ((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!((!env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || ((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[3] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[4] = !((((0 && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || ((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!((0 && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || ((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[5] = !((!(!env_speed_some_high || !(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]))) && adder1_b_invert) || ((!env_speed_some_high || !(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]))) && !(adder1_b_invert)));
    // adder1_b[6] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[7] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[8] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (!env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (!env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[9] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[10] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[11] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && !env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[12] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (!env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (!env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[13] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[14] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[6] && !env_speed_r[5] && !env_speed_r[4] && env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[15] = !(((((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!(((!(!env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[16] = !((((((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (0 && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!((((!env_speed_r[2] && !env_speed_r[1] && env_speed_r[0]) || !((!env_speed_r[2] && env_speed_r[0]) || !env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (0 && env_speed_r[6] && !env_speed_r[5] && env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[17] = !((((!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!((!(!env_speed_r[2] && !env_speed_r[1]) && !env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[18] = !((((((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3])) && adder1_b_invert) || (!((((env_speed_r[2] && !env_speed_r[1] && !env_speed_r[0]) || !(!env_speed_r[1] || !env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && !env_speed_r[4] && env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[19] = !((((env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3])) && adder1_b_invert) || (!((env_speed_r[2] && !(!env_speed_r[1] && !env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && !env_speed_r[3])) && !(adder1_b_invert)));
    // adder1_b[20] = !((env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3] && adder1_b_invert) || (!(env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) && !(adder1_b_invert)));
    
    env_mystery = ((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3]) || (env_speed_r[2] || env_speed_r[1] || env_speed_r[0]));
    adder1_b_invert = env_mystery && env_speed_r[7];

    adder1_b[0] = ~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3] && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[1] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[2] = ~((((~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || ((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~((~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || ((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[3] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[4] = ~((((0 && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || ((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~((0 && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || ((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[5] = ~((~(~(env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) || ~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]))) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || ((~(env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) || ~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]))) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[6] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[7] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[8] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (~env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[9] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[10] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[11] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && ~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[12] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (~env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[13] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[14] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[6] && ~env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[15] = ~(((((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(((~(~env_speed_r[2] || env_speed_r[1]) || env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[16] = ~((((((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (0 && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~((((~env_speed_r[2] && ~env_speed_r[1] && env_speed_r[0]) || ~((~env_speed_r[2] && env_speed_r[0]) || ~env_speed_r[1])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (0 && env_speed_r[6] && ~env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[17] = ~((((~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~((~(~env_speed_r[2] && ~env_speed_r[1]) && ~env_speed_r[0] && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[18] = ~((((((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~((((env_speed_r[2] && ~env_speed_r[1] && ~env_speed_r[0]) || ~(~env_speed_r[1] || ~env_speed_r[0])) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && ~env_speed_r[4] && env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[19] = ~((((env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3])) && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~((env_speed_r[2] && ~(~env_speed_r[1] && ~env_speed_r[0]) && env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) || (env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && ~env_speed_r[3])) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    adder1_b[20] = ~((env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3] && (env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7]) || (~(env_speed_r[6] && env_speed_r[5] && env_speed_r[4] && env_speed_r[3]) && ~((env_speed_r[6] || env_speed_r[5] || env_speed_r[4] || env_speed_r[3] || env_speed_r[2] || env_speed_r[1] || env_speed_r[0]) && env_speed_r[7])));
    // if (adder1_b_invert)
    //   adder1_b = -adder1_b;
    $display("%x", adder1_b);
  end
end

endmodule
