// 79 instances
module cell_LT4 ( // 4-bit Data Latch
  input wire G,
  input wire DA,
  input wire DB,
  input wire DC,
  input wire DD,
  output wire NA,
  output wire PA,
  output wire NB,
  output wire PB,
  output wire NC,
  output wire PC,
  output wire ND,
  output wire PD
);
endmodule

// 3 instances
module cell_DE3 ( // 3:8 Decoder
  input wire B,
  input wire A,
  input wire C,
  output wire X0,
  output wire X1,
  output wire X2,
  output wire X3,
  output wire X4,
  output wire X5,
  output wire X6,
  output wire X7
);
endmodule

// 2 instances
module cell_A2N ( // 2-bit Full Adder
  input wire B2,
  input wire A2,
  input wire B1,
  input wire A1,
  input wire CI,
  output wire CO,
  output wire S2,
  output wire S1
);
endmodule

// 19 instances
module cell_FDQ ( // 4-bit DFF
  input wire CK,
  input wire DA,
  input wire DB,
  input wire DC,
  input wire DD,
  output wire QA,
  output wire QB,
  output wire QC,
  output wire QD
);
endmodule

// 2 instances
module cell_FDR ( // 4-bit DFF with CLEAR
  input wire CL,
  input wire CK,
  input wire DA,
  input wire DB,
  input wire DC,
  input wire DD,
  output wire QA,
  output wire QB,
  output wire QC,
  output wire QD
);
endmodule

// 1 instances
module cell_unkk ( // Unknown K
  input wire A,
  input wire B,
  output wire X
);
endmodule

// 5 instances
module cell_C45 ( // 4-bit Binary Synchronous Up Counter
  input wire DA,
  input wire EN,
  input wire CI,
  input wire CL,
  input wire DB,
  input wire L,
  input wire CK,
  input wire DC,
  input wire DD,
  output wire QA,
  output wire QB,
  output wire CO,
  output wire QC,
  output wire QD
);
endmodule

// 18 instances
module cell_LT2 ( // 1-bit Data Latch
  input wire G,
  input wire D,
  output wire Q,
  output wire XQ
);
endmodule

// 9 instances
module cell_A4H ( // 4-bit Full Adder
  input wire A4,
  input wire B4,
  input wire A3,
  input wire B3,
  input wire A2,
  input wire B2,
  input wire A1,
  input wire B1,
  input wire CI,
  output wire CO,
  output wire S4,
  output wire S3,
  output wire S2,
  output wire S1
);
endmodule

// 13 instances
module cell_FDM ( // DFF
  input wire CK,
  input wire D,
  output wire XQ,
  output wire Q
);
endmodule

// 1 instances
module cell_A1N ( // 1-bit Full Adder
  input wire A,
  input wire B,
  input wire CI,
  output wire CO,
  output wire S
);
endmodule




latch (
  path2452, // INPUT G A104
  R10_D1_IN, // INPUT DA A104
  R10_D0_IN, // INPUT DB A104
  R10_D7_IN, // INPUT DC A104
  R10_D6_IN, // INPUT DD A104
  R10_D5_IN, // INPUT DA A144
  R10_D4_IN, // INPUT DB A144
  R10_D3_IN, // INPUT DC A144
  R10_D2_IN, // INPUT DD A144

  unconnected_A104_NA, // OUTPUT NA A104
  g2511, // OUTPUT PA A104
  unconnected_A104_NB, // OUTPUT NB A104
  g1994, // OUTPUT PB A104
  path2508, // OUTPUT NC A104
  unconnected_A104_PC, // OUTPUT PC A104
  path2507, // OUTPUT ND A104
  unconnected_A104_PD, // OUTPUT PD A104

  path1300, // OUTPUT NA A144
  unconnected_A144_PA, // OUTPUT PA A144
  path2335, // OUTPUT NB A144
  unconnected_A144_PB, // OUTPUT PB A144
  path2336, // OUTPUT NC A144
  unconnected_A144_PC, // OUTPUT PC A144
  unconnected_A144_ND, // OUTPUT ND A144
  g1341, // OUTPUT PD A144
);

latch (
  SYNC_IN, // INPUT G K101
  path1789, // INPUT DA K101
  path1788, // INPUT DB K101
  path1960, // INPUT DC K101
  path1680, // INPUT DD K101
  path1911, // INPUT DA K117
  path2469, // INPUT DB K117
  path2365, // INPUT DC K117
  path1672, // INPUT DD K117
  path1906, // INPUT DA K137
  path1514, // INPUT DB K137
  path1907, // INPUT DC K137
  path2467, // INPUT DD K137
  g2235, // INPUT DA K77
  path1659, // INPUT DB K77
  path2270, // INPUT DC K77
  path2468, // INPUT DD K77
  path1684, // OUTPUT PA K101
  path1683, // OUTPUT PB K101
  path1682, // OUTPUT PC K101
  path1681, // OUTPUT PD K101
  path1912, // OUTPUT PA K117
  path2366, // OUTPUT PB K117
  path2367, // OUTPUT PC K117
  path2368, // OUTPUT PD K117
  path2098, // OUTPUT PA K137
  path1515, // OUTPUT PB K137
  path1517, // OUTPUT PC K137
  path1516, // OUTPUT PD K137
  path1645, // OUTPUT PA K77
  path1656, // OUTPUT PB K77
  path1657, // OUTPUT PC K77
  path1658, // OUTPUT PD K77
);

latch (
  g1731, // INPUT G O80
  g1981, // INPUT DA O80
  g2280, // INPUT DB O80
  g2282, // INPUT DC O80
  g2261, // INPUT DD O80
  g2773, // INPUT DA S77
  path2238, // INPUT DB S77
  path2239, // INPUT DC S77
  path2240, // INPUT DD S77
  g2213, // INPUT DA V123
  g2656, // INPUT DB V123
  g2207, // INPUT DC V123
  g2219, // INPUT DD V123
  g2788, // INPUT DA W103
  g1491, // INPUT DB W103
  g1473, // INPUT DC W103
  path2425, // INPUT DD W103
  path2736, // OUTPUT PA O80
  path1969, // OUTPUT PB O80
  path2316, // OUTPUT PC O80
  path2317, // OUTPUT PD O80
  path2299, // OUTPUT PA S77
  path2298, // OUTPUT PB S77
  path2661, // OUTPUT PC S77
  path2680, // OUTPUT PD S77
  path2644, // OUTPUT PA V123
  path2787, // OUTPUT PB V123
  path2480, // OUTPUT PC V123
  path2635, // OUTPUT PD V123
  path2640, // OUTPUT PA W103
  path2473, // OUTPUT PB W103
  path2660, // OUTPUT PC W103
  path2724, // OUTPUT PD W103
);

latch (
  g1976, // INPUT G O96
  g1981, // INPUT DA O96
  g2280, // INPUT DB O96
  g2282, // INPUT DC O96
  g2261, // INPUT DD O96
  g2773, // INPUT DA S144
  path2238, // INPUT DB S144
  path2239, // INPUT DC S144
  path2240, // INPUT DD S144
  g2213, // INPUT DA V110
  g2656, // INPUT DB V110
  g2207, // INPUT DC V110
  g2219, // INPUT DD V110
  g2788, // INPUT DA W131
  g1491, // INPUT DB W131
  g1473, // INPUT DC W131
  path2425, // INPUT DD W131
  path1968, // OUTPUT PA O96
  path2267, // OUTPUT PB O96
  path2268, // OUTPUT PC O96
  path2262, // OUTPUT PD O96
  path2632, // OUTPUT PA S144
  path2237, // OUTPUT PB S144
  path2305, // OUTPUT PC S144
  path1397, // OUTPUT PD S144
  path2483, // OUTPUT PA V110
  path2641, // OUTPUT PB V110
  path2481, // OUTPUT PC V110
  path2482, // OUTPUT PD V110
  path2723, // OUTPUT PA W131
  path2474, // OUTPUT PB W131
  path2478, // OUTPUT PC W131
  path2472, // OUTPUT PD W131
);

latch (
  r10_ff_clock, // INPUT G P32
  path2403, // INPUT DA P32
  g2256, // INPUT DB P32
  path2180, // INPUT DC P32
  path2406, // INPUT DD P32
  path2763, // INPUT DA H57
  unconnected_H57_DB, // INPUT DB H57
  path2160, // INPUT DC H57
  path2161, // INPUT DD H57
  unconnected_P32_NA, // OUTPUT NA P32
  path2404, // OUTPUT PA P32
  path2734, // OUTPUT NB P32
  path2181, // OUTPUT PB P32
  path2733, // OUTPUT NC P32
  path2735, // OUTPUT PC P32
  path2732, // OUTPUT ND P32
  path2405, // OUTPUT PD P32
  path2708, // OUTPUT NA H57
  path2707, // OUTPUT PA H57
  unconnected_H57_NB, // OUTPUT NB H57
  unconnected_H57_PB, // OUTPUT PB H57
  unconnected_H57_NC, // OUTPUT NC H57
  g1387, // OUTPUT PC H57
  unconnected_H57_ND, // OUTPUT ND H57
  path2512, // OUTPUT PD H57
);

latch (
  g1861, // INPUT G P61
  path1781, // INPUT DA P61
  path1742, // INPUT DB P61
  path2058, // INPUT DC P61
  path1393, // INPUT DD P61
  g1462, // INPUT DA R64
  path1366, // INPUT DB R64
  path1361, // INPUT DC R64
  path2201, // INPUT DD R64
  path1697, // INPUT DA T45
  path1700, // INPUT DB T45
  path2665, // INPUT DC T45
  path1698, // INPUT DD T45
  path1411, // INPUT DA U77
  path1723, // INPUT DB U77
  path1464, // INPUT DC U77
  path1724, // INPUT DD U77
  path1782, // OUTPUT PA P61
  path1741, // OUTPUT PB P61
  path2319, // OUTPUT PC P61
  path1394, // OUTPUT PD P61
  path2408, // OUTPUT PA R64
  path1365, // OUTPUT PB R64
  path1362, // OUTPUT PC R64
  path1729, // OUTPUT PD R64
  path1699, // OUTPUT PA T45
  path2666, // OUTPUT PB T45
  path2242, // OUTPUT PC T45
  path1891, // OUTPUT PD T45
  path1410, // OUTPUT PA U77
  path1465, // OUTPUT PB U77
  path1785, // OUTPUT PC U77
  path1678, // OUTPUT PD U77
);

latch (
  g2048, // INPUT G P80
  g1981, // INPUT DA P80
  g2280, // INPUT DB P80
  g2282, // INPUT DC P80
  g2261, // INPUT DD P80
  g2773, // INPUT DA T90
  path2238, // INPUT DB T90
  path2239, // INPUT DC T90
  path2240, // INPUT DD T90
  g2788, // INPUT DA W116
  g1491, // INPUT DB W116
  g1473, // INPUT DC W116
  path2425, // INPUT DD W116
  g2213, // INPUT DA W77
  g2656, // INPUT DB W77
  g2207, // INPUT DC W77
  g2219, // INPUT DD W77
  path2772, // OUTPUT PA P80
  path2769, // OUTPUT PB P80
  path1939, // OUTPUT PC P80
  path2290, // OUTPUT PD P80
  path1530, // OUTPUT PA T90
  path2751, // OUTPUT PB T90
  path2789, // OUTPUT PC T90
  path2306, // OUTPUT PD T90
  path2284, // OUTPUT PA W116
  path2285, // OUTPUT PB W116
  path1679, // OUTPUT PC W116
  path2645, // OUTPUT PD W116
  path2210, // OUTPUT PA W77
  path2209, // OUTPUT PB W77
  path2216, // OUTPUT PC W77
  path2230, // OUTPUT PD W77
);

latch (
  g1643, // INPUT G Q128
  g1981, // INPUT DA Q128
  g2280, // INPUT DB Q128
  g2282, // INPUT DC Q128
  g2261, // INPUT DD Q128
  g2773, // INPUT DA S131
  path2238, // INPUT DB S131
  path2239, // INPUT DC S131
  path2240, // INPUT DD S131
  g2213, // INPUT DA X144
  g2656, // INPUT DB X144
  g2207, // INPUT DC X144
  g2219, // INPUT DD X144
  g2788, // INPUT DA Y143
  g1491, // INPUT DB Y143
  g1473, // INPUT DC Y143
  path2425, // INPUT DD Y143
  path1973, // OUTPUT PA Q128
  path2770, // OUTPUT PB Q128
  path2273, // OUTPUT PC Q128
  path2276, // OUTPUT PD Q128
  path2303, // OUTPUT PA S131
  path2775, // OUTPUT PB S131
  path2678, // OUTPUT PC S131
  path2677, // OUTPUT PD S131
  path2211, // OUTPUT PA X144
  path2208, // OUTPUT PB X144
  path2217, // OUTPUT PC X144
  path2229, // OUTPUT PD X144
  path1644, // OUTPUT PA Y143
  path1484, // OUTPUT PB Y143
  path2426, // OUTPUT PC Y143
  unconnected_Y143_PD, // OUTPUT PD Y143
);

latch (
  path2231, // INPUT G Q141
  g1981, // INPUT DA Q141
  g2280, // INPUT DB Q141
  g2282, // INPUT DC Q141
  g2261, // INPUT DD Q141
  g2773, // INPUT DA T144
  path2238, // INPUT DB T144
  path2239, // INPUT DC T144
  path2240, // INPUT DD T144
  g2788, // INPUT DA W144
  g1491, // INPUT DB W144
  g1473, // INPUT DC W144
  path2425, // INPUT DD W144
  g2213, // INPUT DA W90
  g2656, // INPUT DB W90
  g2207, // INPUT DC W90
  g2219, // INPUT DD W90
  path2277, // OUTPUT PA Q141
  path2771, // OUTPUT PB Q141
  path2274, // OUTPUT PC Q141
  path2275, // OUTPUT PD Q141
  path2304, // OUTPUT PA T144
  path2294, // OUTPUT PB T144
  path2293, // OUTPUT PC T144
  path1398, // OUTPUT PD T144
  path2648, // OUTPUT PA W144
  path1474, // OUTPUT PB W144
  path2638, // OUTPUT PC W144
  path2228, // OUTPUT PD W144
  path2214, // OUTPUT PA W90
  path2428, // OUTPUT PB W90
  path2427, // OUTPUT PC W90
  path2647, // OUTPUT PD W90
);

latch (
  g2043, // INPUT G R104
  g1981, // INPUT DA R104
  g2280, // INPUT DB R104
  g2282, // INPUT DC R104
  g2261, // INPUT DD R104
  g2773, // INPUT DA S118
  path2238, // INPUT DB S118
  path2239, // INPUT DC S118
  path2240, // INPUT DD S118
  g2213, // INPUT DA X93
  g2656, // INPUT DB X93
  g2207, // INPUT DC X93
  g2219, // INPUT DD X93
  g2788, // INPUT DA Y117
  g1491, // INPUT DB Y117
  g1473, // INPUT DC Y117
  path2425, // INPUT DD Y117
  path2278, // OUTPUT PA R104
  path1971, // OUTPUT PB R104
  path1972, // OUTPUT PC R104
  path2291, // OUTPUT PD R104
  path2750, // OUTPUT PA S118
  path2302, // OUTPUT PB S118
  path2292, // OUTPUT PC S118
  path1904, // OUTPUT PD S118
  path2215, // OUTPUT PA X93
  path2429, // OUTPUT PB X93
  path2430, // OUTPUT PC X93
  path2646, // OUTPUT PD X93
  path2649, // OUTPUT PA Y117
  path2650, // OUTPUT PB Y117
  path2639, // OUTPUT PC Y117
  unconnected_Y117_PD, // OUTPUT PD Y117
);

latch (
  g2436, // INPUT G R77
  g1981, // INPUT DA R77
  g2280, // INPUT DB R77
  g2282, // INPUT DC R77
  g2261, // INPUT DD R77
  g2773, // INPUT DA T131
  path2238, // INPUT DB T131
  path2239, // INPUT DC T131
  path2240, // INPUT DD T131
  g2788, // INPUT DA Y104
  g1491, // INPUT DB Y104
  g1473, // INPUT DC Y104
  path2425, // INPUT DD Y104
  g2213, // INPUT DA Y91
  g2656, // INPUT DB Y91
  g2207, // INPUT DC Y91
  g2219, // INPUT DD Y91
  path2265, // OUTPUT PA R77
  path2266, // OUTPUT PB R77
  path2768, // OUTPUT PC R77
  path2263, // OUTPUT PD R77
  path2631, // OUTPUT PA T131
  path2679, // OUTPUT PB T131
  path2774, // OUTPUT PC T131
  path1903, // OUTPUT PD T131
  path2226, // OUTPUT PA Y104
  path2652, // OUTPUT PB Y104
  path2477, // OUTPUT PC Y104
  path1738, // OUTPUT PD Y104
  path2484, // OUTPUT PA Y91
  path2485, // OUTPUT PB Y91
  path2653, // OUTPUT PC Y91
  path2433, // OUTPUT PD Y91
);

latch (
  g1865, // INPUT G R90
  g1981, // INPUT DA R90
  g2280, // INPUT DB R90
  g2282, // INPUT DC R90
  g2261, // INPUT DD R90
  g2773, // INPUT DA T77
  path2238, // INPUT DB T77
  path2239, // INPUT DC T77
  path2240, // INPUT DD T77
  g2788, // INPUT DA Y130
  g1491, // INPUT DB Y130
  g1473, // INPUT DC Y130
  path2425, // INPUT DD Y130
  g2213, // INPUT DA Y77
  g2656, // INPUT DB Y77
  g2207, // INPUT DC Y77
  g2219, // INPUT DD Y77
  path2264, // OUTPUT PA R90
  path1970, // OUTPUT PB R90
  path2315, // OUTPUT PC R90
  path2314, // OUTPUT PD R90
  path2300, // OUTPUT PA T77
  path2301, // OUTPUT PB T77
  path2295, // OUTPUT PC T77
  path1531, // OUTPUT PD T77
  path2651, // OUTPUT PA Y130
  path2475, // OUTPUT PB Y130
  path2659, // OUTPUT PC Y130
  path2476, // OUTPUT PD Y130
  path2643, // OUTPUT PA Y77
  path2642, // OUTPUT PB Y77
  path2431, // OUTPUT PC Y77
  path2432, // OUTPUT PD Y77
);

latch (
  g2564, // INPUT G B1
  path2576, // INPUT DA B1
  IC19_4_IN, // INPUT DB B1
  g2417, // INPUT DC B1
  IC19_2_IN, // INPUT DD B1
  AG3_IN, // INPUT DA I3
  g1379, // INPUT DB I3
  IC19_6_IN, // INPUT DC I3
  IC19_7_IN, // INPUT DD I3
  path2575, // OUTPUT PA B1
  path2062, // OUTPUT PB B1
  path1374, // OUTPUT PC B1
  path2320, // OUTPUT PD B1
  g1921, // OUTPUT PA I3
  path2112, // OUTPUT PB I3
  path1841, // OUTPUT PC I3
  path1840, // OUTPUT PD I3
);

latch (
  g1750, // INPUT G B104
  g1650, // INPUT DA B104
  g1655, // INPUT DB B104
  g2586, // INPUT DC B104
  g2588, // INPUT DD B104
  g1917, // INPUT DA D104
  g2370, // INPUT DB D104
  g2584, // INPUT DC D104
  g2393, // INPUT DD D104
  g1689, // INPUT DA F77
  g2669, // INPUT DB F77
  g2671, // INPUT DC F77
  g2673, // INPUT DD F77
  g1757, // INPUT DA J127
  path2099, // INPUT DB J127
  g1522, // INPUT DC J127
  g2488, // INPUT DD J127
  path2164, // OUTPUT NA B104
  path2149, // OUTPUT NB B104
  path2148, // OUTPUT NC B104
  path2165, // OUTPUT ND B104
  path2376, // OUTPUT NA D104
  path2063, // OUTPUT NB D104
  path2173, // OUTPUT NC D104
  path2758, // OUTPUT ND D104
  path2741, // OUTPUT NA F77
  path1525, // OUTPUT NB F77
  path1524, // OUTPUT NC F77
  path2399, // OUTPUT ND F77
  path2192, // OUTPUT NA J127
  path1965, // OUTPUT NB J127
  path2762, // OUTPUT NC J127
  path2097, // OUTPUT ND J127
);

latch (
  path1752, // INPUT G B117
  g1650, // INPUT DA B117
  g1655, // INPUT DB B117
  g2586, // INPUT DC B117
  g2588, // INPUT DD B117
  g1917, // INPUT DA D117
  g2370, // INPUT DB D117
  g2584, // INPUT DC D117
  g2393, // INPUT DD D117
  g1689, // INPUT DA F90
  g2669, // INPUT DB F90
  g2671, // INPUT DC F90
  g2673, // INPUT DD F90
  g1757, // INPUT DA J112
  path2099, // INPUT DB J112
  g1522, // INPUT DC J112
  g2488, // INPUT DD J112
  unconnected_B117_NA, // OUTPUT NA B117
  path2754, // OUTPUT NB B117
  path2753, // OUTPUT NC B117
  path2166, // OUTPUT ND B117
  path1615, // OUTPUT NA D117
  path1616, // OUTPUT NB D117
  path2067, // OUTPUT NC D117
  path2066, // OUTPUT ND D117
  path2535, // OUTPUT NA F90
  path2536, // OUTPUT NB F90
  path2103, // OUTPUT NC F90
  path2104, // OUTPUT ND F90
  path1771, // OUTPUT NA J112
  path2504, // OUTPUT NB J112
  path2505, // OUTPUT NC J112
  path2489, // OUTPUT ND J112
);

latch (
  path1607, // INPUT G B130
  g1650, // INPUT DA B130
  g1655, // INPUT DB B130
  g2586, // INPUT DC B130
  g2588, // INPUT DD B130
  g1917, // INPUT DA D131
  g2370, // INPUT DB D131
  g2584, // INPUT DC D131
  g2393, // INPUT DD D131
  g1689, // INPUT DA F142
  g2669, // INPUT DB F142
  g2671, // INPUT DC F142
  g2673, // INPUT DD F142
  g1757, // INPUT DA J140
  path2099, // INPUT DB J140
  g1522, // INPUT DC J140
  g2488, // INPUT DD J140
  path2079, // OUTPUT NA B130
  path2076, // OUTPUT NB B130
  path2089, // OUTPUT NC B130
  path2153, // OUTPUT ND B130
  path1919, // OUTPUT NA D131
  path2064, // OUTPUT NB D131
  path1617, // OUTPUT NC D131
  path2065, // OUTPUT ND D131
  path1610, // OUTPUT NA F142
  path2094, // OUTPUT NB F142
  path2093, // OUTPUT NC F142
  path2397, // OUTPUT ND F142
  path1768, // OUTPUT NA J140
  path1964, // OUTPUT NB J140
  path1769, // OUTPUT NC J140
  path1770, // OUTPUT ND J140
);

latch (
  g1691, // INPUT G B143
  g1650, // INPUT DA B143
  g1655, // INPUT DB B143
  g2586, // INPUT DC B143
  g2588, // INPUT DD B143
  g1917, // INPUT DA D144
  g2370, // INPUT DB D144
  g2584, // INPUT DC D144
  g2393, // INPUT DD D144
  g1689, // INPUT DA F128
  g2669, // INPUT DB F128
  g2671, // INPUT DC F128
  g2673, // INPUT DD F128
  g1757, // INPUT DA H116
  path2099, // INPUT DB H116
  g1522, // INPUT DC H116
  g2488, // INPUT DD H116
  path2078, // OUTPUT NA B143
  path2151, // OUTPUT NB B143
  path2395, // OUTPUT NC B143
  path2396, // OUTPUT ND B143
  path2757, // OUTPUT NA D144
  path2371, // OUTPUT NB D144
  path2374, // OUTPUT NC D144
  path2375, // OUTPUT ND D144
  path2742, // OUTPUT NA F128
  path2102, // OUTPUT NB F128
  path2101, // OUTPUT NC F128
  path1609, // OUTPUT ND F128
  path2193, // OUTPUT NA H116
  path2498, // OUTPUT NB H116
  path1523, // OUTPUT NC H116
  path2497, // OUTPUT ND H116
);

latch (
  path2106, // INPUT G B84
  R10_D1_IN, // INPUT DA B84
  R10_D0_IN, // INPUT DB B84
  unconnected_B84_DC, // INPUT DC B84
  unconnected_B84_DD, // INPUT DD B84
  path2162, // OUTPUT PA B84
  path2740, // OUTPUT PB B84
  unconnected_B84_PC, // OUTPUT PC B84
  unconnected_B84_PD, // OUTPUT PD B84
);

latch (
  g1614, // INPUT G C109
  g1650, // INPUT DA C109
  g1655, // INPUT DB C109
  g2586, // INPUT DC C109
  g2588, // INPUT DD C109
  g1917, // INPUT DA E77
  g2370, // INPUT DB E77
  g2584, // INPUT DC E77
  g2393, // INPUT DD E77
  g1689, // INPUT DA G106
  g2669, // INPUT DB G106
  g2671, // INPUT DC G106
  g2673, // INPUT DD G106
  g1757, // INPUT DA I77
  path2099, // INPUT DB I77
  g1522, // INPUT DC I77
  g2488, // INPUT DD I77
  path2086, // OUTPUT NA C109
  path2087, // OUTPUT NB C109
  path2088, // OUTPUT NC C109
  path2152, // OUTPUT ND C109
  path1918, // OUTPUT NA E77
  path2530, // OUTPUT NB E77
  path2068, // OUTPUT NC E77
  path2069, // OUTPUT ND E77
  path1611, // OUTPUT NA G106
  path2537, // OUTPUT NB G106
  path2092, // OUTPUT NC G106
  path2398, // OUTPUT ND G106
  path2100, // OUTPUT NA I77
  path1758, // OUTPUT NB I77
  path2491, // OUTPUT NC I77
  path2494, // OUTPUT ND I77
);

latch (
  g2156, // INPUT G C144
  g1650, // INPUT DA C144
  g1655, // INPUT DB C144
  g2586, // INPUT DC C144
  g2588, // INPUT DD C144
  g1917, // INPUT DA E90
  g2370, // INPUT DB E90
  g2584, // INPUT DC E90
  g2393, // INPUT DD E90
  g1689, // INPUT DA G143
  g2669, // INPUT DB G143
  g2671, // INPUT DC G143
  g2673, // INPUT DD G143
  g1757, // INPUT DA I90
  path2099, // INPUT DB I90
  g1522, // INPUT DC I90
  g2488, // INPUT DD I90
  path2077, // OUTPUT NA C144
  path2150, // OUTPUT NB C144
  path2394, // OUTPUT NC C144
  path2533, // OUTPUT ND C144
  path2581, // OUTPUT NA E90
  path2372, // OUTPUT NB E90
  path2373, // OUTPUT NC E90
  path2391, // OUTPUT ND E90
  path2157, // OUTPUT NA G143
  path2158, // OUTPUT NB G143
  path2538, // OUTPUT NC G143
  path1608, // OUTPUT ND G143
  path2502, // OUTPUT NA I90
  path2499, // OUTPUT NB I90
  path2500, // OUTPUT NC I90
  path2785, // OUTPUT ND I90
);

latch (
  path2540, // INPUT G C83
  g1650, // INPUT DA C83
  g1655, // INPUT DB C83
  g2586, // INPUT DC C83
  g2588, // INPUT DD C83
  g1917, // INPUT DA D77
  g2370, // INPUT DB D77
  g2584, // INPUT DC D77
  g2393, // INPUT DD D77
  g1689, // INPUT DA G77
  g2669, // INPUT DB G77
  g2671, // INPUT DC G77
  g2673, // INPUT DD G77
  g1757, // INPUT DA H83
  path2099, // INPUT DB H83
  g1522, // INPUT DC H83
  g2488, // INPUT DD H83
  path2163, // OUTPUT NA C83
  path2146, // OUTPUT NB C83
  path2147, // OUTPUT NC C83
  path2755, // OUTPUT ND C83
  path2580, // OUTPUT NA D77
  path2752, // OUTPUT NB D77
  path2389, // OUTPUT NC D77
  path2390, // OUTPUT ND D77
  path2743, // OUTPUT NA G77
  path2159, // OUTPUT NB G77
  path2783, // OUTPUT NC G77
  path2400, // OUTPUT ND G77
  path2490, // OUTPUT NA H83
  path2495, // OUTPUT NB H83
  path2501, // OUTPUT NC H83
  path2096, // OUTPUT ND H83
);

latch (
  path1773, // INPUT G C96
  g1650, // INPUT DA C96
  g1655, // INPUT DB C96
  g2586, // INPUT DC C96
  g2588, // INPUT DD C96
  g1917, // INPUT DA D90
  g2370, // INPUT DB D90
  g2584, // INPUT DC D90
  g2393, // INPUT DD D90
  g1689, // INPUT DA G90
  g2669, // INPUT DB G90
  g2671, // INPUT DC G90
  g2673, // INPUT DD G90
  g1757, // INPUT DA H101
  path2099, // INPUT DB H101
  g1522, // INPUT DC H101
  g2488, // INPUT DD H101
  path2074, // OUTPUT NA C96
  path2075, // OUTPUT NB C96
  path2756, // OUTPUT NC C96
  path2761, // OUTPUT ND C96
  path2760, // OUTPUT NA D90
  path2531, // OUTPUT NB D90
  path2532, // OUTPUT NC D90
  path2759, // OUTPUT ND D90
  path2534, // OUTPUT NA G90
  path2095, // OUTPUT NB G90
  path2539, // OUTPUT NC G90
  path2105, // OUTPUT ND G90
  path1772, // OUTPUT NA H101
  path2496, // OUTPUT NB H101
  path2492, // OUTPUT NC H101
  path2493, // OUTPUT ND H101
);

cell_DE3 L120 ( // 3:8 Decoder
  dac_dec_ia, // INPUT A
  dac_dec_ib, // INPUT B
  dac_dec_ic, // INPUT C
  dac_dec_o0, // OUTPUT X0
  dac_dec_o1, // OUTPUT X1
  dac_dec_o2, // OUTPUT X2
  dac_dec_o3, // OUTPUT X3
  dac_dec_o4, // OUTPUT X4
  dac_dec_o5, // OUTPUT X5
  dac_dec_o6, // OUTPUT X6
  dac_dec_o7, // OUTPUT X7
);

cell_DE3 M103 ( // 3:8 Decoder
  unk_dec_ia, // INPUT A
  unk_dec_ib, // INPUT B
  unk_dec_ic, // INPUT C
  unk_dec_o0, // OUTPUT X0
  unk_dec_o1, // OUTPUT X1
  unk_dec_o2, // OUTPUT X2
  unk_dec_o3, // OUTPUT X3
  unk_dec_o4, // OUTPUT X4
  unk_dec_o5, // OUTPUT X5
  unk_dec_o6, // OUTPUT X6
  unk_dec_o7, // OUTPUT X7
);

cell_DE3 D62 ( // 3:8 Decoder
  cnt_i16_qa, // INPUT A
  cnt_i16_qb, // INPUT B
  cnt_i16_qc, // INPUT C
  cycle_cnt_0, // OUTPUT X0
  cycle_cnt_1, // OUTPUT X1
  cycle_cnt_2, // OUTPUT X2
  cycle_cnt_3, // OUTPUT X3
  cycle_cnt_4, // OUTPUT X4
  cycle_cnt_5, // OUTPUT X5
  cycle_cnt_6, // OUTPUT X6
  cycle_cnt_7, // OUTPUT X7
);

cell_A2N L2 ( // 2-bit Full Adder
  path2421, // INPUT B2
  path2246, // INPUT A2
  path2423, // INPUT B1
  path2692, // INPUT A1
  path2252, // INPUT CI
  path2422, // OUTPUT CO
  path2693, // OUTPUT S2
  path2253, // OUTPUT S1
);

cell_A2N Q61 ( // 2-bit Full Adder
  path2408, // INPUT B2
  path2592, // INPUT A2
  path2408, // INPUT B1
  path2407, // INPUT A1
  path2202, // INPUT CI
  unconnected_Q61_CO, // OUTPUT CO
  path2767, // OUTPUT S2
  path2525, // OUTPUT S1
);

cell_FDQ K50 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  r10_ff_a7, // INPUT DA
  path2420, // INPUT DB
  g2784, // INPUT DC
  path2131, // INPUT DD
  unconnected_K50_QA, // OUTPUT QA
  path2421, // OUTPUT QB
  path2423, // OUTPUT QC
  path2411, // OUTPUT QD
);

cell_FDQ M44 ( // 4-bit DFF
  g1861, // INPUT CK
  path1844, // INPUT DA
  path1845, // INPUT DB
  path2744, // INPUT DC
  unconnected_M44_DD, // INPUT DD
  path2406, // OUTPUT QA
  path2763, // OUTPUT QB
  unconnected_M44_QC, // OUTPUT QC
  unconnected_M44_QD, // OUTPUT QD
);

cell_FDQ M77 ( // 4-bit DFF
  g2564, // INPUT CK
  path2455, // INPUT DA
  path2675, // INPUT DB
  g2446, // INPUT DC
  unconnected_M77_DD, // INPUT DD
  unk_dec_ic, // OUTPUT QA
  unk_dec_ib, // OUTPUT QB
  unk_dec_ia, // OUTPUT QC
  unconnected_M77_QD, // OUTPUT QD
);

cell_FDQ N56 ( // 4-bit DFF
  g1861, // INPUT CK
  unconnected_N56_DA, // INPUT DA
  path1440, // INPUT DB
  path1846, // INPUT DC
  path2254, // INPUT DD
  unconnected_N56_QA, // OUTPUT QA
  path2403, // OUTPUT QB
  g2256, // OUTPUT QC
  path2180, // OUTPUT QD
);

cell_FDQ O117 ( // 4-bit DFF
  g1861, // INPUT CK
  path1848, // INPUT DA
  path2737, // INPUT DB
  path1894, // INPUT DC
  path1893, // INPUT DD
  path1982, // OUTPUT QA
  path2738, // OUTPUT QB
  path1895, // OUTPUT QC
  path1896, // OUTPUT QD
);

cell_FDQ O16 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  AG2_IN, // INPUT DA
  AG1_IN, // INPUT DB
  AG3_IN, // INPUT DC
  ag2_latched, // INPUT DD
  path2776, // OUTPUT QA
  path1833, // OUTPUT QB
  g2034, // OUTPUT QC
  path2602, // OUTPUT QD
);

cell_FDQ O56 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  path2062, // INPUT DA
  path1374, // INPUT DB
  path2320, // INPUT DC
  R6_D1_IN, // INPUT DD
  path2766, // OUTPUT QA
  path1373, // OUTPUT QB
  path2524, // OUTPUT QC
  path2258, // OUTPUT QD
);

cell_FDQ S56 ( // 4-bit DFF
  g1861, // INPUT CK
  path2729, // INPUT DA
  path2686, // INPUT DB
  path2664, // INPUT DC
  path2204, // INPUT DD
  path1890, // OUTPUT QA
  path2629, // OUTPUT QB
  path2663, // OUTPUT QC
  path2662, // OUTPUT QD
);

cell_FDQ T2 ( // 4-bit DFF
  g1861, // INPUT CK
  path2681, // INPUT DA
  path2683, // INPUT DB
  path1887, // INPUT DC
  path1884, // INPUT DD
  path2682, // OUTPUT QA
  path2684, // OUTPUT QB
  path1886, // OUTPUT QC
  path1885, // OUTPUT QD
);

cell_FDQ B16 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  path2321, // INPUT DA
  IC19_4_IN, // INPUT DB
  g2417, // INPUT DC
  IC19_2_IN, // INPUT DD
  path2322, // OUTPUT QA
  path2424, // OUTPUT QB
  path2416, // OUTPUT QC
  path1601, // OUTPUT QD
);

cell_FDQ U56 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  r6_d0_and, // INPUT DA
  R7_D7_IN, // INPUT DB
  R5_D7_IN, // INPUT DC
  r5_d5_and, // INPUT DD
  path2717, // OUTPUT QA
  path2716, // OUTPUT QB
  path2715, // OUTPUT QC
  path2714, // OUTPUT QD
);

cell_FDQ V136 ( // 4-bit DFF
  g1861, // INPUT CK
  path2634, // INPUT DA
  path2633, // INPUT DB
  path1676, // INPUT DC
  path1677, // INPUT DD
  path2479, // OUTPUT QA
  path2636, // OUTPUT QB
  path1675, // OUTPUT QC
  path2637, // OUTPUT QD
);

cell_FDQ X17 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  R6_D2_IN, // INPUT DA
  R7_D2_IN, // INPUT DB
  R7_D1_IN, // INPUT DC
  r5_d1_and, // INPUT DD
  path2018, // OUTPUT QA
  path2572, // OUTPUT QB
  path2711, // OUTPUT QC
  path2521, // OUTPUT QD
);

cell_FDQ X56 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  R5_D2_IN, // INPUT DA
  r5_d6_and, // INPUT DB
  R6_D6_IN, // INPUT DC
  R7_D5_IN, // INPUT DD
  path1421, // OUTPUT QA
  path2616, // OUTPUT QB
  path2712, // OUTPUT QC
  path2624, // OUTPUT QD
);

cell_FDQ Y2 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  r7_d3_and, // INPUT DA
  R5_D0_IN, // INPUT DB
  R6_D4_IN, // INPUT DC
  R7_D4_IN, // INPUT DD
  g2621, // OUTPUT QA
  path1591, // OUTPUT QB
  path2726, // OUTPUT QC
  path2720, // OUTPUT QD
);

cell_FDQ Y35 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  r7_d6_and, // INPUT DA
  R5_D4_IN, // INPUT DB
  R7_D0_IN, // INPUT DC
  r6_d3_and, // INPUT DD
  path2568, // OUTPUT QA
  path1504, // OUTPUT QB
  path2015, // OUTPUT QC
  path2014, // OUTPUT QD
);

cell_FDQ Y56 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  R5_D3_IN, // INPUT DA
  r6_d7_and_2, // INPUT DD
  R6_D5_IN, // INPUT DB
  r6_d7_and, // INPUT DC
  path2727, // OUTPUT QA
  path2713, // OUTPUT QB
  path1450, // OUTPUT QC
  path2625, // OUTPUT QD
);

cell_FDQ E37 ( // 4-bit DFF
  path2702, // INPUT CK
  path2779, // INPUT DA
  path2780, // INPUT DB
  path2781, // INPUT DC
  unconnected_E37_DD, // INPUT DD
  path2703, // OUTPUT QA
  path2704, // OUTPUT QB
  path2705, // OUTPUT QC
  unconnected_E37_QD, // OUTPUT QD
);

cell_FDQ J1 ( // 4-bit DFF
  cycle_odd_inv, // INPUT CK
  path2112, // INPUT DA
  path1841, // INPUT DB
  path1840, // INPUT DC
  path2575, // INPUT DD
  path2113, // OUTPUT QA
  path1839, // OUTPUT QB
  path2574, // OUTPUT QC
  path1842, // OUTPUT QD
);

cell_FDR A117 ( // 4-bit DFF with CLEAR
  MPX1_IOM, // INPUT CL
  MPX1_IN, // INPUT CK
  R10_D7_IN, // INPUT DA
  R10_D6_IN, // INPUT DB
  R10_D5_IN, // INPUT DC
  R10_D4_IN, // INPUT DD
  r10_ff_a117_d7, // OUTPUT QA
  r10_ff_a117_d6, // OUTPUT QB
  r10_ff_a117_d5, // OUTPUT QC
  r10_ff_a117_d4, // OUTPUT QD
);
cell_FDR A77 ( // 4-bit DFF with CLEAR
  MPX1_IOM, // INPUT CL
  MPX1_IN, // INPUT CK
  R10_D3_IN, // INPUT DA
  R10_D2_IN, // INPUT DB
  R10_D1_IN, // INPUT DC
  R10_D0_IN, // INPUT DD
  r10_ff_a77_d3, // OUTPUT QA
  r10_ff_a77_d2, // OUTPUT QB
  r10_ff_a77_d1, // OUTPUT QC
  r10_ff_a77_d0, // OUTPUT QD
);

cell_unkk C58 ( // Unknown K
  path2695, // INPUT A
  path2544, // INPUT B
  g1691, // OUTPUT X
);

cell_C45 C1 ( // 4-bit Binary Synchronous Up Counter
  unconnected_C1_EN, // INPUT EN
  path1986, // INPUT CL
  unconnected_C1_L, // INPUT L
  r10_ff_clock, // INPUT CK
  unconnected_C1_CI, // INPUT CI
  
  unconnected_C1_DA, // INPUT DA
  unconnected_C1_DB, // INPUT DB
  g2136, // INPUT DC
  unconnected_C1_DD, // INPUT DD
  
  path2696, // OUTPUT QA
  unconnected_C1_QB, // OUTPUT QB
  unconnected_C1_QC, // OUTPUT QC
  path1984, // OUTPUT QD
  
  unconnected_C1_CO, // OUTPUT CO
);

cell_C45 D1 ( // 4-bit Binary Synchronous Up Counter
  path2108, // INPUT EN
  path2323, // INPUT CL
  unconnected_D1_L, // INPUT L
  r10_ff_clock, // INPUT CK
  unconnected_D1_CI, // INPUT CI
  
  unconnected_D1_DA, // INPUT DA
  unconnected_D1_DB, // INPUT DB
  g2136, // INPUT DC
  unconnected_D1_DD, // INPUT DD
  
  g107, // OUTPUT QA
  path1987, // OUTPUT QB
  path2362, // OUTPUT QC
  g2361, // OUTPUT QD
  
  unconnected_D1_CO, // OUTPUT CO
);

cell_C45 G29 ( // 4-bit Binary Synchronous Up Counter
  r10_ff_a5, // INPUT EN
  FSYNC_IN, // INPUT CL
  path1791, // INPUT L
  r10_ff_clock, // INPUT CK
  unconnected_G29_CI, // INPUT CI
  
  path1715, // INPUT DA
  g2782, // INPUT DB
  g1994, // INPUT DC
  unconnected_G29_DD, // INPUT DD
  
  g1720, // OUTPUT QA
  g2446, // OUTPUT QB
  path2675, // OUTPUT QC
  path2455, // OUTPUT QD
  
  clock_low_sr, // OUTPUT CO
);

cell_C45 H1 ( // 4-bit Binary Synchronous Up Counter
  path1988, // INPUT EN
  FSYNC_IN, // INPUT CL
  unconnected_H1_L, // INPUT L
  r10_ff_clock, // INPUT CK
  unconnected_H1_CI, // INPUT CI
  
  unconnected_H1_DA, // INPUT DA
  unconnected_H1_DB, // INPUT DB
  g2136, // INPUT DC
  unconnected_H1_DD, // INPUT DD
  
  MPX1_OUT, // OUTPUT QA
  unconnected_H1_QB, // OUTPUT QB
  path2780, // OUTPUT QC
  path2781, // OUTPUT QD
  
  path2109, // OUTPUT CO
);

cell_C45 I16 ( // 4-bit Binary Synchronous Up Counter
  unconnected_I16_EN, // INPUT EN
  FSYNC_IN, // INPUT CL
  unconnected_I16_L, // INPUT L
  SYNC_IN, // INPUT CK
  g2698, // INPUT CI
  
  unconnected_I16_DA, // INPUT DA
  unconnected_I16_DB, // INPUT DB
  path2744, // INPUT DC
  path2675, // INPUT DD
  
  cnt_i16_qa, // OUTPUT QA
  cnt_i16_qb, // OUTPUT QB
  cnt_i16_qc, // OUTPUT QC
  cnt_i16_qd, // OUTPUT QD
  
  unconnected_I16_CO, // OUTPUT CO
);

cell_LT2 N109 ( // 1-bit Data Latch
  g2043, // INPUT G
  path2035, // INPUT D
  path2233, // OUTPUT Q
  unconnected_N109_XQ, // OUTPUT XQ
);

cell_LT2 N113 ( // 1-bit Data Latch
  path2231, // INPUT G
  path2035, // INPUT D
  path2232, // OUTPUT Q
  unconnected_N113_XQ, // OUTPUT XQ
);

cell_LT2 N122 ( // 1-bit Data Latch
  g1643, // INPUT G
  path2035, // INPUT D
  path2764, // OUTPUT Q
  unconnected_N122_XQ, // OUTPUT XQ
);

cell_LT2 N126 ( // 1-bit Data Latch
  g1976, // INPUT G
  path2035, // INPUT D
  path2223, // OUTPUT Q
  unconnected_N126_XQ, // OUTPUT XQ
);

cell_LT2 N77 ( // 1-bit Data Latch
  g2436, // INPUT G
  path2035, // INPUT D
  path2222, // OUTPUT Q
  unconnected_N77_XQ, // OUTPUT XQ
);

cell_LT2 N81 ( // 1-bit Data Latch
  g1865, // INPUT G
  path2035, // INPUT D
  path1866, // OUTPUT Q
  unconnected_N81_XQ, // OUTPUT XQ
);

cell_LT2 N85 ( // 1-bit Data Latch
  g1731, // INPUT G
  path2035, // INPUT D
  path1867, // OUTPUT Q
  unconnected_N85_XQ, // OUTPUT XQ
);

cell_LT2 N89 ( // 1-bit Data Latch
  g2048, // INPUT G
  path2035, // INPUT D
  path2765, // OUTPUT Q
  unconnected_N89_XQ, // OUTPUT XQ
);

cell_LT2 O5 ( // 1-bit Data Latch
  g2564, // INPUT G
  AG2_IN, // INPUT D
  ag2_latched, // OUTPUT Q
  unconnected_O5_XQ, // OUTPUT XQ
);

cell_LT2 O9 ( // 1-bit Data Latch
  g2564, // INPUT G
  AG1_IN, // INPUT D
  ag1_latched, // OUTPUT Q
  unconnected_O9_XQ, // OUTPUT XQ
);

cell_LT2 R117 ( // 1-bit Data Latch
  g2048, // INPUT G
  path2055, // INPUT D
  path2049, // OUTPUT Q
  unconnected_R117_XQ, // OUTPUT XQ
);

cell_LT2 R121 ( // 1-bit Data Latch
  g1731, // INPUT G
  path2055, // INPUT D
  path2050, // OUTPUT Q
  unconnected_R121_XQ, // OUTPUT XQ
);

cell_LT2 R137 ( // 1-bit Data Latch
  g1865, // INPUT G
  path2055, // INPUT D
  path1528, // OUTPUT Q
  unconnected_R137_XQ, // OUTPUT XQ
);

cell_LT2 R141 ( // 1-bit Data Latch
  g2043, // INPUT G
  path2055, // INPUT D
  path2052, // OUTPUT Q
  unconnected_R141_XQ, // OUTPUT XQ
);

cell_LT2 R145 ( // 1-bit Data Latch
  g1643, // INPUT G
  path2055, // INPUT D
  path2051, // OUTPUT Q
  unconnected_R145_XQ, // OUTPUT XQ
);

cell_LT2 R149 ( // 1-bit Data Latch
  g1976, // INPUT G
  path2055, // INPUT D
  path2054, // OUTPUT Q
  unconnected_R149_XQ, // OUTPUT XQ
);

cell_LT2 R153 ( // 1-bit Data Latch
  path2231, // INPUT G
  path2055, // INPUT D
  path2053, // OUTPUT Q
  unconnected_R153_XQ, // OUTPUT XQ
);

cell_LT2 S102 ( // 1-bit Data Latch
  g2436, // INPUT G
  path2055, // INPUT D
  path1529, // OUTPUT Q
  unconnected_S102_XQ, // OUTPUT XQ
);

cell_A4H L27 ( // 4-bit Full Adder
  path2411, // INPUT A4
  path2410, // INPUT B4
  path2322, // INPUT A3
  path2249, // INPUT B3
  path2424, // INPUT A2
  path2412, // INPUT B2
  path2416, // INPUT A1
  path2415, // INPUT B1
  path2137, // INPUT CI
  path2252, // OUTPUT CO
  path2251, // OUTPUT S4
  path2250, // OUTPUT S3
  r10_ff_a10, // OUTPUT S2
  r10_ff_a9, // OUTPUT S1
);

cell_A4H N5 ( // 4-bit Full Adder
  path1842, // INPUT A4
  path1843, // INPUT B4
  path2766, // INPUT A3
  path2566, // INPUT B3
  path1373, // INPUT A2
  path1372, // INPUT B2
  path2524, // INPUT A1
  path1414, // INPUT B1
  g2562, // INPUT CI
  path2590, // OUTPUT CO
  r10_ff_a4, // OUTPUT S4
  r10_ff_a3, // OUTPUT S3
  r10_ff_a2, // OUTPUT S2
  r10_ff_a7, // OUTPUT S1
);

cell_A4H P98 ( // 4-bit Full Adder
  path1891, // INPUT A4
  path1892, // INPUT B4
  path1782, // INPUT A3
  path1783, // INPUT B3
  path1741, // INPUT A2
  path1740, // INPUT B2
  path2319, // INPUT A1
  path2318, // INPUT B1
  path1509, // INPUT CI
  path1883, // OUTPUT CO
  path1848, // OUTPUT S4
  path2737, // OUTPUT S3
  path1894, // OUTPUT S2
  path1893, // OUTPUT S1
);

cell_A4H R4 ( // 4-bit Full Adder
  path2408, // INPUT A4
  path2409, // INPUT B4
  path2408, // INPUT A3
  path2730, // INPUT B3
  path1365, // INPUT A2
  path1364, // INPUT B2
  path1362, // INPUT A1
  path1363, // INPUT B1
  path2203, // INPUT CI
  path2202, // OUTPUT CO
  path2729, // OUTPUT S4
  path2686, // OUTPUT S3
  path2664, // OUTPUT S2
  path2204, // OUTPUT S1
);

cell_A4H S3 ( // 4-bit Full Adder
  path1729, // INPUT A4
  path1728, // INPUT B4
  path1699, // INPUT A3
  path2243, // INPUT B3
  path2666, // INPUT A2
  path2728, // INPUT B2
  path2242, // INPUT A1
  path2241, // INPUT B1
  path1883, // INPUT CI
  path2203, // OUTPUT CO
  path2681, // OUTPUT S4
  path2683, // OUTPUT S3
  path1887, // OUTPUT S2
  path1884, // OUTPUT S1
);

cell_A4H U107 ( // 4-bit Full Adder
  path1394, // INPUT A4
  path2307, // INPUT B4
  path1410, // INPUT A3
  path1409, // INPUT B3
  path1465, // INPUT A2
  path1466, // INPUT B2
  path1785, // INPUT A1
  path1784, // INPUT B1
  path1678, // INPUT CI
  path1509, // OUTPUT CO
  path2634, // OUTPUT S4
  path2633, // OUTPUT S3
  path1676, // OUTPUT S2
  path1677, // OUTPUT S1
);

cell_A4H V4 ( // 4-bit Full Adder
  path2603, // INPUT A4
  path1504, // INPUT B4
  path2614, // INPUT A3
  path2015, // INPUT B3
  path2013, // INPUT A2
  path2014, // INPUT B2
  path1420, // INPUT A1
  path1421, // INPUT B1
  path1997, // INPUT CI
  path1597, // OUTPUT CO
  path2604, // OUTPUT S4
  path2749, // OUTPUT S3
  path1598, // OUTPUT S2
  path2017, // OUTPUT S1
);

cell_A4H W1 ( // 4-bit Full Adder
  path2009, // INPUT A4
  path2616, // INPUT B4
  path2571, // INPUT A3
  path2712, // INPUT B3
  path2786, // INPUT A2
  path2624, // INPUT B2
  path2622, // INPUT A1
  path2625, // INPUT B1
  unconnected_W1_CI, // INPUT CI
  path1997, // OUTPUT CO
  path2615, // OUTPUT S4
  path2016, // OUTPUT S3
  path2520, // OUTPUT S2
  path2626, // OUTPUT S1
);

cell_A4H J27 ( // 4-bit Full Adder
  path1601, // INPUT A4
  path1600, // INPUT B4
  path2113, // INPUT A3
  path2523, // INPUT B3
  path1839, // INPUT A2
  path2573, // INPUT B2
  path2574, // INPUT A1
  path2709, // INPUT B1
  path2590, // INPUT CI
  path2137, // OUTPUT CO
  r10_ff_a8, // OUTPUT S4
  r10_ff_a7, // OUTPUT S3
  r10_ff_a6, // OUTPUT S2
  r10_ff_a5, // OUTPUT S1
);

cell_FDM A2 ( // DFF
  r10_ff_clock, // INPUT CK
  r10_ff_a10, // INPUT D
  unconnected_A2_XQ, // OUTPUT XQ
  R10_A10_OUT, // OUTPUT Q
);

cell_FDM A17 ( // DFF
  path1330, // INPUT CK
  path1328, // INPUT D
  unconnected_A17_XQ, // OUTPUT XQ
  path1329, // OUTPUT Q
);

cell_FDM A23 ( // DFF
  r10_ff_clock, // INPUT CK
  r10_ff_a8, // INPUT D
  unconnected_A23_XQ, // OUTPUT XQ
  R10_A8_OUT, // OUTPUT Q
);

cell_FDM A29 ( // DFF
  r10_ff_clock, // INPUT CK
  r10_ff_a5, // INPUT D
  unconnected_A29_XQ, // OUTPUT XQ
  R10_A5_OUT, // OUTPUT Q
);

cell_FDM A45 ( // DFF
  r10_ff_clock, // INPUT CK
  r10_ff_a4, // INPUT D
  unconnected_A45_XQ, // OUTPUT XQ
  R10_A4_OUT, // OUTPUT Q
);

cell_FDM A51 ( // DFF
  r10_ff_clock, // INPUT CK
  r10_ff_a7, // INPUT D
  unconnected_A51_XQ, // OUTPUT XQ
  R10_A1_OUT, // OUTPUT Q
);

cell_FDM A71 ( // DFF
  r10_ff_clock, // INPUT CK
  r10_ff_a7, // INPUT D
  unconnected_A71_XQ, // OUTPUT XQ
  R10_A7_OUT, // OUTPUT Q
);

cell_FDM P51 ( // DFF
  path2184, // INPUT CK
  path2767, // INPUT D
  path2591, // OUTPUT XQ
  unconnected_P51_Q, // OUTPUT Q
);

cell_FDM Q42 ( // DFF
  path2184, // INPUT CK
  path2525, // INPUT D
  path2056, // OUTPUT XQ
  unconnected_Q42_Q, // OUTPUT Q
);

cell_FDM B77 ( // DFF
  r10_ff_clock, // INPUT CK
  r10_ff_a3, // INPUT D
  unconnected_B77_XQ, // OUTPUT XQ
  R10_A3_OUT, // OUTPUT Q
);

cell_FDM B98 ( // DFF
  r10_ff_clock, // INPUT CK
  r10_ff_a6, // INPUT D
  unconnected_B98_XQ, // OUTPUT XQ
  R10_A6_OUT, // OUTPUT Q
);

cell_FDM C77 ( // DFF
  r10_ff_clock, // INPUT CK
  r10_ff_a2, // INPUT D
  unconnected_C77_XQ, // OUTPUT XQ
  R10_A2_OUT, // OUTPUT Q
);

cell_FDM E116 ( // DFF
  r10_ff_clock, // INPUT CK
  r10_ff_a9, // INPUT D
  unconnected_E116_XQ, // OUTPUT XQ
  R10_A9_OUT, // OUTPUT Q
);

cell_A1N V69 ( // 1-bit Full Adder
  path2002, // INPUT A
  path2568, // INPUT B
  path1597, // INPUT CI
  path2605, // OUTPUT CO
  path1596, // OUTPUT S
);

assign cycle0_n = cycle_cnt_0 || SYNC_IN || ~cnt_i16_qd;
assign cycle1_n = cycle_cnt_1 || SYNC_IN || ~cnt_i16_qd;
assign cycle2_n = cycle_cnt_2 || SYNC_IN || ~cnt_i16_qd;
assign cycle3_n = cycle_cnt_3 || SYNC_IN || ~cnt_i16_qd;
assign cycle4_n = cycle_cnt_4 || SYNC_IN || ~cnt_i16_qd;
assign cycle5_n = cycle_cnt_5 || SYNC_IN || ~cnt_i16_qd;
assign cycle6_n = cycle_cnt_6 || SYNC_IN || ~cnt_i16_qd;
assign cycle7_n = cycle_cnt_7 || SYNC_IN || ~cnt_i16_qd;
assign cycle8_p = cycle_cnt_0 || SYNC_IN || cnt_i16_qd;
assign cycle9_p = cycle_cnt_1 || SYNC_IN || cnt_i16_qd;
assign cycle10_p = cycle_cnt_2 || SYNC_IN || cnt_i16_qd;
assign cycle11_p = cycle_cnt_3 || SYNC_IN || cnt_i16_qd;
assign cycle12_p = cycle_cnt_4 || SYNC_IN || cnt_i16_qd;
assign cycle13_p = cycle_cnt_5 || SYNC_IN || cnt_i16_qd;
assign cycle14_p = cycle_cnt_6 || SYNC_IN || cnt_i16_qd;
assign cycle15_p = cycle_cnt_7 || SYNC_IN || cnt_i16_qd;

assign cycle_odd = cycle7_n && cycle5_n && cycle3_n && cycle1_n && cycle15_p && cycle13_p && cycle11_p && cycle9_p;
assign cycle_even = cycle6_n && cycle4_n && cycle2_n && cycle0_n && cycle14_p && cycle12_p && cycle10_p && cycle8_p;
assign cycle_odd_or_even = ~cycle_odd || ~cycle_even;
assign cycle_odd_inv = ~cycle_odd;

assign tmp1 = (path1984 && path2696 && SR_SEL_IN) || (clock_low_sr && ~SR_SEL_IN);

assign DAC1_OUT = ~(~(~(((~SR_SEL_IN && g107) || path1987 || path2362 || g2361) && (MPX1_OUT || path2779 || path2780 || path2781)) && r10_ff_a77_d2) && ~(~((path2375 && ~dac_dec_o0) || (path2391 && ~dac_dec_o1) || (path2758 && ~dac_dec_o2) || (path2390 && ~dac_dec_o3) || (path2066 && ~dac_dec_o4) || (path2759 && ~dac_dec_o5) || (path2065 && ~dac_dec_o6) || (path2069 && ~dac_dec_o7)) && ~r10_ff_a77_d2));
assign DAC2_OUT = ~(~((~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0) && r10_ff_a77_d2) && ~(~((path2374 && ~dac_dec_o0) || (path2373 && ~dac_dec_o1) || (path2173 && ~dac_dec_o2) || (path2389 && ~dac_dec_o3) || (path2067 && ~dac_dec_o4) || (path2532 && ~dac_dec_o5) || (path1617 && ~dac_dec_o6) || (path2068 && ~dac_dec_o7)) && ~r10_ff_a77_d2));
assign DAC3_OUT = ~(~(~((path2645 && path2455 && ~path2675 && g2446) || (path2225 && path2455 && ~path2675 && ~g2446) || (path2228 && ~path2455 && path2675 && g2446) || (path2227 && ~path2455 && path2675 && ~g2446) || (path2724 && ~path2455 && ~path2675 && g2446) || (path2476 && ~path2455 && ~path2675 && ~g2446) || (path2472 && path2455 && path2675 && g2446) || (path1738 && path2455 && path2675 && ~g2446)) && r10_ff_a77_d2) && ~(~((path2371 && ~dac_dec_o0) || (path2372 && ~dac_dec_o1) || (path2063 && ~dac_dec_o2) || (path2752 && ~dac_dec_o3) || (path1616 && ~dac_dec_o4) || (path2531 && ~dac_dec_o5) || (path2064 && ~dac_dec_o6) || (path2530 && ~dac_dec_o7)) && ~r10_ff_a77_d2));
assign DAC4_OUT = ~(~(~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && r10_ff_a77_d2) && ~(~((path2757 && ~dac_dec_o0) || (path2581 && ~dac_dec_o1) || (path2376 && ~dac_dec_o2) || (path2580 && ~dac_dec_o3) || (path1615 && ~dac_dec_o4) || (path2760 && ~dac_dec_o5) || (path1919 && ~dac_dec_o6) || (path1918 && ~dac_dec_o7)) && ~r10_ff_a77_d2));
assign DAC5_OUT = ~(~(path2763 && r10_ff_a77_d2) && ~(~((path2497 && ~dac_dec_o0) || (path2785 && ~dac_dec_o1) || (path2097 && ~dac_dec_o2) || (path2096 && ~dac_dec_o3) || (path2489 && ~dac_dec_o4) || (path2493 && ~dac_dec_o5) || (path1770 && ~dac_dec_o6) || (path2494 && ~dac_dec_o7)) && ~r10_ff_a77_d2));
assign DAC6_OUT = ~(~(path2406 && r10_ff_a77_d2) && ~(~((path1523 && ~dac_dec_o0) || (path2500 && ~dac_dec_o1) || (path2762 && ~dac_dec_o2) || (path2501 && ~dac_dec_o3) || (path2505 && ~dac_dec_o4) || (path2492 && ~dac_dec_o5) || (path1769 && ~dac_dec_o6) || (path2491 && ~dac_dec_o7)) && ~r10_ff_a77_d2));
assign DAC7_OUT = ~(~(path2180 && r10_ff_a77_d2) && ~(~((path2498 && ~dac_dec_o0) || (path2499 && ~dac_dec_o1) || (path1965 && ~dac_dec_o2) || (path2495 && ~dac_dec_o3) || (path2504 && ~dac_dec_o4) || (path2496 && ~dac_dec_o5) || (path1964 && ~dac_dec_o6) || (path1758 && ~dac_dec_o7)) && ~r10_ff_a77_d2));
assign DAC8_OUT = ~(~(g2256 && r10_ff_a77_d2) && ~(~((path2193 && ~dac_dec_o0) || (path2502 && ~dac_dec_o1) || (path2192 && ~dac_dec_o2) || (path2490 && ~dac_dec_o3) || (path1771 && ~dac_dec_o4) || (path1772 && ~dac_dec_o5) || (path1768 && ~dac_dec_o6) || (path2100 && ~dac_dec_o7)) && ~r10_ff_a77_d2));
assign DAC9_OUT = ~(~(path2403 && r10_ff_a77_d2) && ~(~((path1609 && ~dac_dec_o0) || (path1608 && ~dac_dec_o1) || (path2399 && ~dac_dec_o2) || (path2400 && ~dac_dec_o3) || (path2104 && ~dac_dec_o4) || (path2105 && ~dac_dec_o5) || (path2397 && ~dac_dec_o6) || (path2398 && ~dac_dec_o7)) && ~r10_ff_a77_d2));
assign DAC10_OUT = ~((path2101 && ~dac_dec_o0) || (path2538 && ~dac_dec_o1) || (path1524 && ~dac_dec_o2) || (path2783 && ~dac_dec_o3) || (path2103 && ~dac_dec_o4) || (path2539 && ~dac_dec_o5) || (path2093 && ~dac_dec_o6) || (path2092 && ~dac_dec_o7));
assign DAC11_OUT = ~((path2102 && ~dac_dec_o0) || (path2158 && ~dac_dec_o1) || (path1525 && ~dac_dec_o2) || (path2159 && ~dac_dec_o3) || (path2536 && ~dac_dec_o4) || (path2095 && ~dac_dec_o5) || (path2094 && ~dac_dec_o6) || (path2537 && ~dac_dec_o7));
assign DAC12_OUT = ~((path2742 && ~dac_dec_o0) || (path2157 && ~dac_dec_o1) || (path2741 && ~dac_dec_o2) || (path2743 && ~dac_dec_o3) || (path2535 && ~dac_dec_o4) || (path2534 && ~dac_dec_o5) || (path1610 && ~dac_dec_o6) || (path1611 && ~dac_dec_o7));
assign DAC13_OUT = ~((path2396 && ~dac_dec_o0) || (path2533 && ~dac_dec_o1) || (path2165 && ~dac_dec_o2) || (path2755 && ~dac_dec_o3) || (path2166 && ~dac_dec_o4) || (path2761 && ~dac_dec_o5) || (path2153 && ~dac_dec_o6) || (path2152 && ~dac_dec_o7));
assign DAC14_OUT = ~((path2395 && ~dac_dec_o0) || (path2394 && ~dac_dec_o1) || (path2148 && ~dac_dec_o2) || (path2147 && ~dac_dec_o3) || (path2753 && ~dac_dec_o4) || (path2756 && ~dac_dec_o5) || (path2089 && ~dac_dec_o6) || (path2088 && ~dac_dec_o7));
assign DAC15_OUT = ~((path2151 && ~dac_dec_o0) || (path2150 && ~dac_dec_o1) || (path2149 && ~dac_dec_o2) || (path2146 && ~dac_dec_o3) || (path2754 && ~dac_dec_o4) || (path2075 && ~dac_dec_o5) || (path2076 && ~dac_dec_o6) || (path2087 && ~dac_dec_o7));
assign DAC16_OUT = (path2078 && ~dac_dec_o0) || (path2077 && ~dac_dec_o1) || (path2164 && ~dac_dec_o2) || (path2163 && ~dac_dec_o3) || (unconnected_C133_E1 && ~dac_dec_o4) || (path2074 && ~dac_dec_o5) || (path2079 && ~dac_dec_o6) || (path2086 && ~dac_dec_o7);

assign FSYNC_OUT = ~(path2109 && g2361 && g107 && (tmp1 || r10_ff_a117_d4));
assign MPX2_OUT = ~((((~((path2645 && path2455 && ~path2675 && g2446) || (path2225 && path2455 && ~path2675 && ~g2446) || (path2228 && ~path2455 && path2675 && g2446) || (path2227 && ~path2455 && path2675 && ~g2446) || (path2724 && ~path2455 && ~path2675 && g2446) || (path2476 && ~path2455 && ~path2675 && ~g2446) || (path2472 && path2455 && path2675 && g2446) || (path1738 && path2455 && path2675 && ~g2446)) && ~cycle_odd_or_even) || (cycle_odd_or_even && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)))) && r10_ff_a117_d7) || (MPX1_OUT && ~r10_ff_a117_d7));
assign R10_A0_OUT = cycle_odd_or_even;

assign r10_ff_clock = ~cycle_odd_or_even;
assign dac_dec_ia = (r10_ff_a77_d1 && g2446) || (~r10_ff_a77_d1 && path2703);
assign dac_dec_ib = (r10_ff_a77_d1 && path2675) || (~r10_ff_a77_d1 && path2704);
assign dac_dec_ic = (r10_ff_a77_d1 && path2455) || (~r10_ff_a77_d1 && path2705);

assign r5_d1_and = ~((~R5_D1_IN && r10_ff_a117_d5) || (R5_D1_IN && ~r10_ff_a117_d5));
assign r5_d5_and = ~((~R5_D5_IN && r10_ff_a117_d5) || (R5_D5_IN && ~r10_ff_a117_d5));
assign r5_d6_and = ~((~R5_D6_IN && r10_ff_a117_d5) || (R5_D6_IN && ~r10_ff_a117_d5));
assign r6_d0_and = ~((~R6_D0_IN && r10_ff_a117_d5) || (R6_D0_IN && ~r10_ff_a117_d5));
assign r6_d3_and = ~((~R6_D3_IN && r10_ff_a117_d5) || (R6_D3_IN && ~r10_ff_a117_d5));
assign r6_d7_and = ~((R6_D7_IN && ~r10_ff_a117_d5) || ~(R6_D7_IN || ~r10_ff_a117_d5) || g1921);
assign r6_d7_and_2 = ~((R6_D7_IN && ~r10_ff_a117_d5) || ~(R6_D7_IN || ~r10_ff_a117_d5) || ~g1921);
assign r7_d3_and = ~((~R7_D3_IN && r10_ff_a117_d5) || (R7_D3_IN && ~r10_ff_a117_d5));
assign r7_d6_and = ~((~R7_D6_IN && r10_ff_a117_d5) || (R7_D6_IN && ~r10_ff_a117_d5));

assign g1865 = unk_dec_o0 || cycle_odd_or_even;
assign g1731 = unk_dec_o1 || cycle_odd_or_even;
assign g2043 = unk_dec_o2 || cycle_odd_or_even;
assign path2231 = unk_dec_o3 || cycle_odd_or_even;
assign g1643 = unk_dec_o4 || cycle_odd_or_even;
assign g2048 = unk_dec_o5 || cycle_odd_or_even;
assign g2436 = unk_dec_o6 || cycle_odd_or_even;
assign g1976 = unk_dec_o7 || cycle_odd_or_even;

assign g1379 = ~((~IC19_1_IN && r10_ff_a117_d5) || (IC19_1_IN && ~r10_ff_a117_d5));
assign g1462 = path2404;
assign g1473 = path1675;
assign g1491 = path2636;
assign g1522 = ~path1517;
assign g1614 = ~(~(cycle3_n || ~r10_ff_a77_d3) || ~(cycle2_n || ~(r10_ff_a77_d3 || path1329)));
assign g1650 = ~path1645;
assign g1655 = ~path1656;
assign g1689 = ~path1684;
assign g1750 = ~(~(cycle9_p || ~r10_ff_a77_d3) || ~(cycle8_p || ~(r10_ff_a77_d3 || path1329)));
assign g1757 = ~path2098;
assign g1861 = cycle_odd_or_even;
assign g1917 = ~path1912;
assign g1981 = path1982;
assign g2136 = SYNC_IN || cnt_i16_qd;
assign g2156 = ~(~(cycle7_n || ~r10_ff_a77_d3) || ~(cycle6_n || ~(r10_ff_a77_d3 || path1329)));
assign g2207 = path1886;
assign g2213 = path2682;
assign g2219 = path1885;
assign g2235 = ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446));
assign g2261 = path1896;
assign g2280 = path2738;
assign g2282 = path1895;
assign g2370 = ~path2366;
assign g2393 = ~path2368;
assign g2417 = ~((~IC19_3_IN && r10_ff_a117_d5) || (IC19_3_IN && ~r10_ff_a117_d5));
assign g2488 = ~path1516;
assign g2562 = ~((~path1300 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~path2507 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (~path2508 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (unconnected_D49_D1 && ~path2181 && ~path2735 && ~path2732 && ~path2708));
assign g2564 = cycle_even;
assign g2584 = ~path2367;
assign g2586 = ~path1657;
assign g2588 = ~path1658;
assign g2656 = path2684;
assign g2669 = ~path1683;
assign g2671 = ~path1682;
assign g2673 = ~path1681;
assign g2698 = SYNC_IN || ~cnt_i16_qd;
assign g2773 = path1890;
assign g2782 = ~(g2361 && g107 && ~(~tmp1 && ~r10_ff_a117_d4));
assign g2784 = IC19_6_IN || ag1_latched;
assign g2788 = path2479;
assign path1328 = ~(((~SR_SEL_IN && g107) || path1987 || path2362 || g2361) && (MPX1_OUT || path2779 || path2780 || path2781));
assign path1330 = ~cycle3_n;
assign path1361 = ~((((~path2508 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~path2181 && ~path2735 && ~path2405 && ~path2708)) && path2404) || (~((~path2508 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~path2181 && ~path2735 && ~path2405 && ~path2708)) && ~path2404));
assign path1363 = ~(~((path2306 && path2455 && ~path2675 && g2446) || (path2677 && path2455 && ~path2675 && ~g2446) || (path1398 && ~path2455 && path2675 && g2446) || (path1904 && ~path2455 && path2675 && ~g2446) || (path2680 && ~path2455 && ~path2675 && g2446) || (path1531 && ~path2455 && ~path2675 && ~g2446) || (path1397 && path2455 && path2675 && g2446) || (path1903 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path1364 = ~(~((path2789 && path2455 && ~path2675 && g2446) || (path2678 && path2455 && ~path2675 && ~g2446) || (path2293 && ~path2455 && path2675 && g2446) || (path2292 && ~path2455 && path2675 && ~g2446) || (path2661 && ~path2455 && ~path2675 && g2446) || (path2295 && ~path2455 && ~path2675 && ~g2446) || (path2305 && path2455 && path2675 && g2446) || (path2774 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path1366 = ~((~(~path2181 && ~path2735 && ~path2405 && ~path2707) && ~path2404) || (~path2181 && ~path2735 && ~path2405 && ~path2707 && path2404));
assign path1372 = ~(~(path2713 && ~g1720) && ~(unconnected_T23_A1 && g1720));
assign path1393 = ~((~((path2512 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (g1387 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (g1994 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g2511 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g1341 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (~path2336 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2335 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path1300 && ~path2181 && ~path2733 && ~path2732 && ~path2708)) && ~((~path2507 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path2508 && ~path2734 && ~path2735 && ~path2405 && ~path2708) || (~path2734 && ~path2735 && ~path2732 && ~path2707)) && ~path2404) || (~(~((path2512 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (g1387 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (g1994 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g2511 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g1341 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (~path2336 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2335 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path1300 && ~path2181 && ~path2733 && ~path2732 && ~path2708)) && ~((~path2507 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path2508 && ~path2734 && ~path2735 && ~path2405 && ~path2708) || (~path2734 && ~path2735 && ~path2732 && ~path2707))) && path2404));
assign path1409 = ~(~((path2285 && path2455 && ~path2675 && g2446) || (path1484 && path2455 && ~path2675 && ~g2446) || (path1474 && ~path2455 && path2675 && g2446) || (path2650 && ~path2455 && path2675 && ~g2446) || (path2473 && ~path2455 && ~path2675 && g2446) || (path2475 && ~path2455 && ~path2675 && ~g2446) || (path2474 && path2455 && path2675 && g2446) || (path2652 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path1411 = ~((~((path2512 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (g1387 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g1994 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g2511 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g1341 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2336 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2335 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path1300 && ~path2734 && ~path2735 && ~path2405 && ~path2707)) && ~((~path2507 && ~path2734 && ~path2735 && ~path2405 && ~path2708) || (~path2508 && ~path2734 && ~path2735 && ~path2732 && ~path2707) || (~path2734 && ~path2735 && ~path2732 && ~path2708)) && ~path2404) || (~(~((path2512 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (g1387 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g1994 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g2511 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g1341 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2336 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2335 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path1300 && ~path2734 && ~path2735 && ~path2405 && ~path2707)) && ~((~path2507 && ~path2734 && ~path2735 && ~path2405 && ~path2708) || (~path2508 && ~path2734 && ~path2735 && ~path2732 && ~path2707) || (~path2734 && ~path2735 && ~path2732 && ~path2708))) && path2404));
assign path1414 = ~(~(path1450 && ~g1720) && ~(unconnected_T75_A1 && g1720));
assign path1420 = ~(~(~path2776 && path1833 && ~g2034 && path2602) && ~(path2776 && ~unconnected_O49_A && ~g2034 && path2602) && ~(path2776 && ~unconnected_O49_A && g2034 && ~path2602) && ~(path2776 && ~unconnected_O49_A && g2034 && path2602));
assign path1440 = ~(~(g2621 && ~g1720) && ~(path2258 && g1720));
assign path1464 = ~((~((path2512 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g1387 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g1994 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (g2511 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (g1341 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path2336 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path2335 && ~path2734 && ~path2735 && ~path2405 && ~path2708) || (~path1300 && ~path2734 && ~path2735 && ~path2732 && ~path2707)) && ~((~path2507 && ~path2734 && ~path2735 && ~path2732 && ~path2708) || (~path2508 && ~path2734 && ~path2733 && ~path2405 && ~path2707) || (~path2734 && ~path2733 && ~path2405 && ~path2708)) && ~path2404) || (~(~((path2512 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g1387 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g1994 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (g2511 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (g1341 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path2336 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path2335 && ~path2734 && ~path2735 && ~path2405 && ~path2708) || (~path1300 && ~path2734 && ~path2735 && ~path2732 && ~path2707)) && ~((~path2507 && ~path2734 && ~path2735 && ~path2732 && ~path2708) || (~path2508 && ~path2734 && ~path2733 && ~path2405 && ~path2707) || (~path2734 && ~path2733 && ~path2405 && ~path2708))) && path2404));
assign path1466 = ~(~((path1679 && path2455 && ~path2675 && g2446) || (path2426 && path2455 && ~path2675 && ~g2446) || (path2638 && ~path2455 && path2675 && g2446) || (path2639 && ~path2455 && path2675 && ~g2446) || (path2660 && ~path2455 && ~path2675 && g2446) || (path2659 && ~path2455 && ~path2675 && ~g2446) || (path2478 && path2455 && path2675 && g2446) || (path2477 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path1514 = ~(~(~((path2772 && path2455 && ~path2675 && g2446) || (path1973 && path2455 && ~path2675 && ~g2446) || (path2277 && ~path2455 && path2675 && g2446) || (path2278 && ~path2455 && path2675 && ~g2446) || (path2736 && ~path2455 && ~path2675 && g2446) || (path2264 && ~path2455 && ~path2675 && ~g2446) || (path1968 && path2455 && path2675 && g2446) || (path2265 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path1600 = ~(~(path2714 && ~g1720) && ~(path2016 && g1720));
assign path1607 = ~(~(cycle1_n || ~r10_ff_a77_d3) || ~(cycle0_n || ~(r10_ff_a77_d3 || path1329)));
assign path1659 = ~(~(~((path1530 && path2455 && ~path2675 && g2446) || (path2303 && path2455 && ~path2675 && ~g2446) || (path2304 && ~path2455 && path2675 && g2446) || (path2750 && ~path2455 && path2675 && ~g2446) || (path2299 && ~path2455 && ~path2675 && g2446) || (path2300 && ~path2455 && ~path2675 && ~g2446) || (path2632 && path2455 && path2675 && g2446) || (path2631 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path1672 = ~(~(~((path1679 && path2455 && ~path2675 && g2446) || (path2426 && path2455 && ~path2675 && ~g2446) || (path2638 && ~path2455 && path2675 && g2446) || (path2639 && ~path2455 && path2675 && ~g2446) || (path2660 && ~path2455 && ~path2675 && g2446) || (path2659 && ~path2455 && ~path2675 && ~g2446) || (path2478 && path2455 && path2675 && g2446) || (path2477 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path1680 = ~(~(~((path2216 && path2455 && ~path2675 && g2446) || (path2217 && path2455 && ~path2675 && ~g2446) || (path2427 && ~path2455 && path2675 && g2446) || (path2430 && ~path2455 && path2675 && ~g2446) || (path2480 && ~path2455 && ~path2675 && g2446) || (path2431 && ~path2455 && ~path2675 && ~g2446) || (path2481 && path2455 && path2675 && g2446) || (path2653 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path1697 = ~((((~path1300 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~path2507 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (~path2508 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (unconnected_D49_D1 && ~path2181 && ~path2735 && ~path2732 && ~path2708)) && path2404) || (~((~path1300 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~path2507 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (~path2508 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (unconnected_D49_D1 && ~path2181 && ~path2735 && ~path2732 && ~path2708)) && ~path2404));
assign path1698 = ~((((unconnected_F1_A1 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2508 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2507 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (~path1300 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (~path2335 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (~path2336 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (g1341 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~((~IC19_1_IN && r10_ff_a117_d5) || (IC19_1_IN && ~r10_ff_a117_d5)) && unconnected_F1_H2)) && path2404) || (~((unconnected_F1_A1 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2508 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2507 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (~path1300 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (~path2335 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (~path2336 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (g1341 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~((~IC19_1_IN && r10_ff_a117_d5) || (IC19_1_IN && ~r10_ff_a117_d5)) && unconnected_F1_H2)) && ~path2404));
assign path1700 = ~((~((~path2508 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (~path2507 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (~path1300 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (~path2335 && ~path2181 && ~path2735 && ~path2405 && ~path2707)) && ~(~path2181 && ~path2733 && ~path2405 && ~path2707) && ~path2404) || (~(~((~path2508 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (~path2507 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (~path1300 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (~path2335 && ~path2181 && ~path2735 && ~path2405 && ~path2707)) && ~(~path2181 && ~path2733 && ~path2405 && ~path2707)) && path2404));
assign path1715 = ~g1720;
assign path1723 = ~((~((path2512 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g1387 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g1994 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g2511 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (g1341 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2336 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path2335 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path1300 && ~path2734 && ~path2735 && ~path2405 && ~path2708)) && ~((~path2507 && ~path2734 && ~path2735 && ~path2732 && ~path2707) || (~path2508 && ~path2734 && ~path2735 && ~path2732 && ~path2708) || (~path2734 && ~path2733 && ~path2405 && ~path2707)) && ~path2404) || (~(~((path2512 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g1387 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g1994 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g2511 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (g1341 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2336 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path2335 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path1300 && ~path2734 && ~path2735 && ~path2405 && ~path2708)) && ~((~path2507 && ~path2734 && ~path2735 && ~path2732 && ~path2707) || (~path2508 && ~path2734 && ~path2735 && ~path2732 && ~path2708) || (~path2734 && ~path2733 && ~path2405 && ~path2707))) && path2404));
assign path1724 = ~((~((path2512 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g1387 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (g1994 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (g2511 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (g1341 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path2336 && ~path2734 && ~path2735 && ~path2405 && ~path2708) || (~path2335 && ~path2734 && ~path2735 && ~path2732 && ~path2707) || (~path1300 && ~path2734 && ~path2735 && ~path2732 && ~path2708)) && ~((~path2507 && ~path2734 && ~path2733 && ~path2405 && ~path2707) || (~path2508 && ~path2734 && ~path2733 && ~path2405 && ~path2708) || (~path2734 && ~path2733 && ~path2732 && ~path2707)) && ~path2404) || (~(~((path2512 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g1387 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (g1994 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (g2511 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (g1341 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path2336 && ~path2734 && ~path2735 && ~path2405 && ~path2708) || (~path2335 && ~path2734 && ~path2735 && ~path2732 && ~path2707) || (~path1300 && ~path2734 && ~path2735 && ~path2732 && ~path2708)) && ~((~path2507 && ~path2734 && ~path2733 && ~path2405 && ~path2707) || (~path2508 && ~path2734 && ~path2733 && ~path2405 && ~path2708) || (~path2734 && ~path2733 && ~path2732 && ~path2707))) && path2404));
assign path1728 = ~(~((path2210 && path2455 && ~path2675 && g2446) || (path2211 && path2455 && ~path2675 && ~g2446) || (path2214 && ~path2455 && path2675 && g2446) || (path2215 && ~path2455 && path2675 && ~g2446) || (path2644 && ~path2455 && ~path2675 && g2446) || (path2643 && ~path2455 && ~path2675 && ~g2446) || (path2483 && path2455 && path2675 && g2446) || (path2484 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path1740 = ~(~((path1939 && path2455 && ~path2675 && g2446) || (path2273 && path2455 && ~path2675 && ~g2446) || (path2274 && ~path2455 && path2675 && g2446) || (path1972 && ~path2455 && path2675 && ~g2446) || (path2316 && ~path2455 && ~path2675 && g2446) || (path2315 && ~path2455 && ~path2675 && ~g2446) || (path2268 && path2455 && path2675 && g2446) || (path2768 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path1742 = ~((~((path2779 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path2508 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path2507 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path1300 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2335 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (~path2336 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g1341 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g2511 && ~path2181 && ~path2735 && ~path2405 && ~path2708)) && ~(g1994 && ~path2181 && ~path2735 && ~path2405 && ~path2707) && ~path2404) || (~(~((path2779 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path2508 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path2507 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path1300 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2335 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (~path2336 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g1341 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g2511 && ~path2181 && ~path2735 && ~path2405 && ~path2708)) && ~(g1994 && ~path2181 && ~path2735 && ~path2405 && ~path2707)) && path2404));
assign path1752 = ~(~(cycle13_p || ~r10_ff_a77_d3) || ~(cycle12_p || ~(r10_ff_a77_d3 || path1329)));
assign path1773 = ~(~(cycle15_p || ~r10_ff_a77_d3) || ~(cycle14_p || ~(r10_ff_a77_d3 || path1329)));
assign path1781 = ~((((~cycle_odd_or_even && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path2508 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2507 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path1300 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (~path2335 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (~path2336 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g1341 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (g2511 && ~path2181 && ~path2735 && ~path2405 && ~path2707)) && path2404) || (~((~cycle_odd_or_even && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path2508 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2507 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path1300 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (~path2335 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (~path2336 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g1341 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (g2511 && ~path2181 && ~path2735 && ~path2405 && ~path2707)) && ~path2404));
assign path1783 = ~(~((path2769 && path2455 && ~path2675 && g2446) || (path2770 && path2455 && ~path2675 && ~g2446) || (path2771 && ~path2455 && path2675 && g2446) || (path1971 && ~path2455 && path2675 && ~g2446) || (path1969 && ~path2455 && ~path2675 && g2446) || (path1970 && ~path2455 && ~path2675 && ~g2446) || (path2267 && path2455 && path2675 && g2446) || (path2266 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path1784 = ~(~((path2645 && path2455 && ~path2675 && g2446) || (path2225 && path2455 && ~path2675 && ~g2446) || (path2228 && ~path2455 && path2675 && g2446) || (path2227 && ~path2455 && path2675 && ~g2446) || (path2724 && ~path2455 && ~path2675 && g2446) || (path2476 && ~path2455 && ~path2675 && ~g2446) || (path2472 && path2455 && path2675 && g2446) || (path1738 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path1788 = ~(~(~((path2210 && path2455 && ~path2675 && g2446) || (path2211 && path2455 && ~path2675 && ~g2446) || (path2214 && ~path2455 && path2675 && g2446) || (path2215 && ~path2455 && path2675 && ~g2446) || (path2644 && ~path2455 && ~path2675 && g2446) || (path2643 && ~path2455 && ~path2675 && ~g2446) || (path2483 && path2455 && path2675 && g2446) || (path2484 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path1789 = ~(~(~((path2306 && path2455 && ~path2675 && g2446) || (path2677 && path2455 && ~path2675 && ~g2446) || (path1398 && ~path2455 && path2675 && g2446) || (path1904 && ~path2455 && path2675 && ~g2446) || (path2680 && ~path2455 && ~path2675 && g2446) || (path1531 && ~path2455 && ~path2675 && ~g2446) || (path1397 && path2455 && path2675 && g2446) || (path1903 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path1791 = ~r10_ff_a117_d6;
assign path1843 = ~(~(path2521 && ~g1720) && ~(unconnected_U12_A1 && g1720));
assign path1844 = path2251 || path2422;
assign path1845 = path2250 || path2422;
assign path1846 = path2693 || path2422;
assign path1892 = ~(~((path2772 && path2455 && ~path2675 && g2446) || (path1973 && path2455 && ~path2675 && ~g2446) || (path2277 && ~path2455 && path2675 && g2446) || (path2278 && ~path2455 && path2675 && ~g2446) || (path2736 && ~path2455 && ~path2675 && g2446) || (path2264 && ~path2455 && ~path2675 && ~g2446) || (path1968 && path2455 && path2675 && g2446) || (path2265 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path1906 = ~(~(~((path2230 && path2455 && ~path2675 && g2446) || (path2229 && path2455 && ~path2675 && ~g2446) || (path2647 && ~path2455 && path2675 && g2446) || (path2646 && ~path2455 && path2675 && ~g2446) || (path2635 && ~path2455 && ~path2675 && g2446) || (path2432 && ~path2455 && ~path2675 && ~g2446) || (path2482 && path2455 && path2675 && g2446) || (path2433 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path1907 = ~(~(~((path2769 && path2455 && ~path2675 && g2446) || (path2770 && path2455 && ~path2675 && ~g2446) || (path2771 && ~path2455 && path2675 && g2446) || (path1971 && ~path2455 && path2675 && ~g2446) || (path1969 && ~path2455 && ~path2675 && g2446) || (path1970 && ~path2455 && ~path2675 && ~g2446) || (path2267 && path2455 && path2675 && g2446) || (path2266 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path1911 = ~(~(~((path2290 && path2455 && ~path2675 && g2446) || (path2276 && path2455 && ~path2675 && ~g2446) || (path2275 && ~path2455 && path2675 && g2446) || (path2291 && ~path2455 && path2675 && ~g2446) || (path2317 && ~path2455 && ~path2675 && g2446) || (path2314 && ~path2455 && ~path2675 && ~g2446) || (path2262 && path2455 && path2675 && g2446) || (path2263 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path1960 = ~(~(~((path2209 && path2455 && ~path2675 && g2446) || (path2208 && path2455 && ~path2675 && ~g2446) || (path2428 && ~path2455 && path2675 && g2446) || (path2429 && ~path2455 && path2675 && ~g2446) || (path2787 && ~path2455 && ~path2675 && g2446) || (path2642 && ~path2455 && ~path2675 && ~g2446) || (path2641 && path2455 && path2675 && g2446) || (path2485 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path1986 = FSYNC_IN && ~(path1984 && path2696);
assign path1988 = g2361 && g107 && ~(~tmp1 && ~r10_ff_a117_d4);
assign path2002 = ~path2776 && ~unconnected_O49_A && ~g2034 && ~path2602;
assign path2009 = ~(unconnected_X5_A1 && ~(~path2776 && ~unconnected_O49_A && g2034 && path2602) && ~(~path2776 && path1833 && g2034 && ~path2602) && ~(path2776 && ~unconnected_O49_A && ~g2034 && path2602) && ~(path2776 && path1833 && ~g2034 && ~path2602) && ~(path2776 && path1833 && ~g2034 && path2602));
assign path2013 = ~(~(~path2776 && ~unconnected_O49_A && ~g2034 && ~path2602) && ~(~path2776 && ~unconnected_O49_A && g2034 && ~path2602) && ~(~path2776 && path1833 && ~g2034 && path2602) && ~(~path2776 && path1833 && g2034 && ~path2602) && ~(~path2776 && path1833 && g2034 && path2602) && ~(path2776 && ~unconnected_O49_A && ~g2034 && ~path2602));
assign path2035 = ~path2591;
assign path2055 = ~path2056;
assign path2058 = ~((~((~path2508 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path2507 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path1300 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2335 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2336 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g1341 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g2511 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g1994 && ~path2181 && ~path2735 && ~path2405 && ~path2708)) && ~((g1387 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~path2734 && ~path2735 && ~path2405 && ~path2708)) && ~path2404) || (~(~((~path2508 && ~path2734 && ~path2735 && ~path2405 && ~path2707) || (~path2507 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path1300 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2335 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2336 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g1341 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g2511 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g1994 && ~path2181 && ~path2735 && ~path2405 && ~path2708)) && ~((g1387 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~path2734 && ~path2735 && ~path2405 && ~path2708))) && path2404));
assign path2099 = ~path1515;
assign path2106 = ~(~cycle_odd_or_even && unconnected_J101_A2);
assign path2108 = ~(~tmp1 && ~r10_ff_a117_d4);
assign path2131 = IC19_7_IN || ag1_latched;
assign path2160 = path2162;
assign path2161 = path2740;
assign path2184 = ~cycle_odd_or_even;
assign path2201 = ~((((~path2507 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~path2508 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (~path2181 && ~path2735 && ~path2732 && ~path2707)) && path2404) || (~((~path2507 && ~path2181 && ~path2735 && ~path2405 && ~path2707) || (~path2508 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (~path2181 && ~path2735 && ~path2732 && ~path2707)) && ~path2404));
assign path2238 = path2629;
assign path2239 = path2663;
assign path2240 = path2662;
assign path2241 = ~(~((path2230 && path2455 && ~path2675 && g2446) || (path2229 && path2455 && ~path2675 && ~g2446) || (path2647 && ~path2455 && path2675 && g2446) || (path2646 && ~path2455 && path2675 && ~g2446) || (path2635 && ~path2455 && ~path2675 && g2446) || (path2432 && ~path2455 && ~path2675 && ~g2446) || (path2482 && path2455 && path2675 && g2446) || (path2433 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path2243 = ~(~((path2209 && path2455 && ~path2675 && g2446) || (path2208 && path2455 && ~path2675 && ~g2446) || (path2428 && ~path2455 && path2675 && g2446) || (path2429 && ~path2455 && path2675 && ~g2446) || (path2787 && ~path2455 && ~path2675 && g2446) || (path2642 && ~path2455 && ~path2675 && ~g2446) || (path2641 && path2455 && path2675 && g2446) || (path2485 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path2246 = ~(~(path1591 && ~g1720) && ~((path1596 || path2605) && g1720));
assign path2249 = ~(~(path2717 && ~g1720) && ~((path1598 || path2605) && g1720));
assign path2254 = path2253 || path2422;
assign path2270 = ~(~(~((path2751 && path2455 && ~path2675 && g2446) || (path2775 && path2455 && ~path2675 && ~g2446) || (path2294 && ~path2455 && path2675 && g2446) || (path2302 && ~path2455 && path2675 && ~g2446) || (path2298 && ~path2455 && ~path2675 && g2446) || (path2301 && ~path2455 && ~path2675 && ~g2446) || (path2237 && path2455 && path2675 && g2446) || (path2679 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path2307 = ~(~((path2284 && path2455 && ~path2675 && g2446) || (path1644 && path2455 && ~path2675 && ~g2446) || (path2648 && ~path2455 && path2675 && g2446) || (path2649 && ~path2455 && path2675 && ~g2446) || (path2640 && ~path2455 && ~path2675 && g2446) || (path2651 && ~path2455 && ~path2675 && ~g2446) || (path2723 && path2455 && path2675 && g2446) || (path2226 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path2318 = ~(~((path2290 && path2455 && ~path2675 && g2446) || (path2276 && path2455 && ~path2675 && ~g2446) || (path2275 && ~path2455 && path2675 && g2446) || (path2291 && ~path2455 && path2675 && ~g2446) || (path2317 && ~path2455 && ~path2675 && g2446) || (path2314 && ~path2455 && ~path2675 && ~g2446) || (path2262 && path2455 && path2675 && g2446) || (path2263 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path2321 = ~((~IC19_5_IN && r10_ff_a117_d5) || (IC19_5_IN && ~r10_ff_a117_d5)) || ag1_latched;
assign path2323 = FSYNC_IN && ~(g2361 && g107 && ~(~tmp1 && ~r10_ff_a117_d4));
assign path2365 = ~(~(~((path2285 && path2455 && ~path2675 && g2446) || (path1484 && path2455 && ~path2675 && ~g2446) || (path1474 && ~path2455 && path2675 && g2446) || (path2650 && ~path2455 && path2675 && ~g2446) || (path2473 && ~path2455 && ~path2675 && g2446) || (path2475 && ~path2455 && ~path2675 && ~g2446) || (path2474 && path2455 && path2675 && g2446) || (path2652 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path2407 = ~(~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path2409 = ~(~((path1530 && path2455 && ~path2675 && g2446) || (path2303 && path2455 && ~path2675 && ~g2446) || (path2304 && ~path2455 && path2675 && g2446) || (path2750 && ~path2455 && path2675 && ~g2446) || (path2299 && ~path2455 && ~path2675 && g2446) || (path2300 && ~path2455 && ~path2675 && ~g2446) || (path2632 && path2455 && path2675 && g2446) || (path2631 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path2410 = ~(~(path2720 && ~g1720) && ~((path2749 || path2605) && g1720));
assign path2412 = ~(~(path2716 && ~g1720) && ~(path2017 && g1720));
assign path2415 = ~(~(path2715 && ~g1720) && ~(path2615 && g1720));
assign path2420 = ~((~IC19_1_IN && r10_ff_a117_d5) || (IC19_1_IN && ~r10_ff_a117_d5)) || ag1_latched;
assign path2425 = path2637;
assign path2452 = ~cycle_odd_or_even && unconnected_J101_A2;
assign path2467 = ~(~(~((path1939 && path2455 && ~path2675 && g2446) || (path2273 && path2455 && ~path2675 && ~g2446) || (path2274 && ~path2455 && path2675 && g2446) || (path1972 && ~path2455 && path2675 && ~g2446) || (path2316 && ~path2455 && ~path2675 && g2446) || (path2315 && ~path2455 && ~path2675 && ~g2446) || (path2268 && path2455 && path2675 && g2446) || (path2768 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path2468 = ~(~(~((path2789 && path2455 && ~path2675 && g2446) || (path2678 && path2455 && ~path2675 && ~g2446) || (path2293 && ~path2455 && path2675 && g2446) || (path2292 && ~path2455 && path2675 && ~g2446) || (path2661 && ~path2455 && ~path2675 && g2446) || (path2295 && ~path2455 && ~path2675 && ~g2446) || (path2305 && path2455 && path2675 && g2446) || (path2774 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path2469 = ~(~(~((path2284 && path2455 && ~path2675 && g2446) || (path1644 && path2455 && ~path2675 && ~g2446) || (path2648 && ~path2455 && path2675 && g2446) || (path2649 && ~path2455 && path2675 && ~g2446) || (path2640 && ~path2455 && ~path2675 && g2446) || (path2651 && ~path2455 && ~path2675 && ~g2446) || (path2723 && path2455 && path2675 && g2446) || (path2226 && path2455 && path2675 && ~g2446)) || (((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7)) || (((path2049 && path2455 && ~path2675 && g2446) || (path2051 && path2455 && ~path2675 && ~g2446) || (path2053 && ~path2455 && path2675 && g2446) || (path2052 && ~path2455 && path2675 && ~g2446) || (path2050 && ~path2455 && ~path2675 && g2446) || (path1528 && ~path2455 && ~path2675 && ~g2446) || (path2054 && path2455 && path2675 && g2446) || (path1529 && path2455 && path2675 && ~g2446)) && ~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) && ~r10_ff_a117_d7));
assign path2523 = ~(~(path2018 && ~g1720) && ~(path2520 && g1720));
assign path2540 = ~(~(cycle11_p || ~r10_ff_a77_d3) || ~(cycle10_p || ~(r10_ff_a77_d3 || path1329)));
assign path2544 = ~(cycle4_n || ~(r10_ff_a77_d3 || path1329));
assign path2566 = ~(~(path2727 && ~g1720) && ~(unconnected_U14_A1 && g1720));
assign path2571 = ~(g2621 && ~(~path2776 && ~unconnected_O49_A && g2034 && path2602) && ~(~path2776 && path1833 && ~g2034 && path2602) && ~(~path2776 && path1833 && g2034 && ~path2602) && ~(~path2776 && path1833 && g2034 && path2602) && ~(path2776 && ~unconnected_O49_A && g2034 && ~path2602) && ~(path2776 && path1833 && ~g2034 && ~path2602) && ~(path2776 && path1833 && g2034 && ~path2602));
assign path2573 = ~(~(path2572 && ~g1720) && ~(path2626 && g1720));
assign path2576 = ~((~IC19_5_IN && r10_ff_a117_d5) || (IC19_5_IN && ~r10_ff_a117_d5));
assign path2592 = ~(~((path2765 && path2455 && ~path2675 && g2446) || (path2764 && path2455 && ~path2675 && ~g2446) || (path2232 && ~path2455 && path2675 && g2446) || (path2233 && ~path2455 && path2675 && ~g2446) || (path1867 && ~path2455 && ~path2675 && g2446) || (path1866 && ~path2455 && ~path2675 && ~g2446) || (path2223 && path2455 && path2675 && g2446) || (path2222 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path2603 = ~(~(~path2776 && ~unconnected_O49_A && ~g2034 && ~path2602) && ~(~path2776 && ~unconnected_O49_A && ~g2034 && path2602));
assign path2614 = ~(~(~path2776 && ~unconnected_O49_A && ~g2034 && ~path2602) && ~(~path2776 && ~unconnected_O49_A && g2034 && ~path2602) && ~(~path2776 && ~unconnected_O49_A && g2034 && path2602) && ~(~path2776 && path1833 && ~g2034 && ~path2602));
assign path2622 = ~(~(~path2776 && ~unconnected_O49_A && g2034 && path2602) && ~(~path2776 && path1833 && g2034 && ~path2602) && ~(path2776 && ~unconnected_O49_A && ~g2034 && path2602) && ~(path2776 && ~unconnected_O49_A && g2034 && path2602) && ~(path2776 && path1833 && ~g2034 && ~path2602) && ~(path2776 && path1833 && g2034 && path2602));
assign path2665 = ~((((unconnected_F12_A1 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2508 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (~path2507 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (~path1300 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (~path2335 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (~path2336 && ~path2181 && ~path2735 && ~path2405 && ~path2707)) && path2404) || (~((unconnected_F12_A1 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2508 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (~path2507 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (~path1300 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (~path2335 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (~path2336 && ~path2181 && ~path2735 && ~path2405 && ~path2707)) && ~path2404));
assign path2692 = ~(~(path2726 && ~g1720) && ~((path2604 || path2605) && g1720));
assign path2695 = ~(cycle5_n || ~r10_ff_a77_d3);
assign path2702 = cycle7_n;
assign path2709 = ~(~(path2711 && ~g1720) && ~(unconnected_U46_A1 && g1720));
assign path2728 = ~(~((path2216 && path2455 && ~path2675 && g2446) || (path2217 && path2455 && ~path2675 && ~g2446) || (path2427 && ~path2455 && path2675 && g2446) || (path2430 && ~path2455 && path2675 && ~g2446) || (path2480 && ~path2455 && ~path2675 && g2446) || (path2431 && ~path2455 && ~path2675 && ~g2446) || (path2481 && path2455 && path2675 && g2446) || (path2653 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path2730 = ~(~((path2751 && path2455 && ~path2675 && g2446) || (path2775 && path2455 && ~path2675 && ~g2446) || (path2294 && ~path2455 && path2675 && g2446) || (path2302 && ~path2455 && path2675 && ~g2446) || (path2298 && ~path2455 && ~path2675 && g2446) || (path2301 && ~path2455 && ~path2675 && ~g2446) || (path2237 && path2455 && path2675 && g2446) || (path2679 && path2455 && path2675 && ~g2446)) || ~(~(r10_ff_a77_d3 || path1329) || g1720) || r10_ff_a77_d0);
assign path2744 = ~(~((path2512 && ~path2181 && ~path2735 && ~path2405 && ~path2708) || (g1387 && ~path2181 && ~path2735 && ~path2732 && ~path2707) || (g1994 && ~path2181 && ~path2735 && ~path2732 && ~path2708) || (g2511 && ~path2181 && ~path2733 && ~path2405 && ~path2707) || (g1341 && ~path2181 && ~path2733 && ~path2405 && ~path2708) || (~path2336 && ~path2181 && ~path2733 && ~path2732 && ~path2707) || (~path2335 && ~path2181 && ~path2733 && ~path2732 && ~path2708) || (~path1300 && ~path2734 && ~path2735 && ~path2405 && ~path2707)) && ~((~path2507 && ~path2734 && ~path2735 && ~path2405 && ~path2708) || (~path2508 && ~path2734 && ~path2735 && ~path2732 && ~path2707) || (~path2734 && ~path2735 && ~path2732 && ~path2708)));
assign path2786 = ~(unconnected_X50_A1 && ~(~path2776 && path1833 && ~g2034 && path2602) && ~(~path2776 && path1833 && g2034 && path2602) && ~(path2776 && ~unconnected_O49_A && ~g2034 && path2602) && ~(path2776 && ~unconnected_O49_A && g2034 && ~path2602) && ~(path2776 && path1833 && ~g2034 && path2602) && ~(path2776 && path1833 && g2034 && ~path2602) && ~(path2776 && path1833 && g2034 && path2602));
